module rtu_rob (
    clk,
    rst_clk,
    y_rtu_rob_stall_ctrl,
    idu_rtu_rob_iid_req_vld,
    idu_rtu_rob_create_vld,
    idu_rtu_rob_create_opcode,
    idu_rtu_rob_create_funct3,
    idu_rtu_rob_create_pc,
    idu_rtu_rob_create_src1,
    idu_rtu_rob_create_src1_vld,
    idu_rtu_rob_create_psrc1,
    idu_rtu_rob_create_src2,
    idu_rtu_rob_create_src2_vld,
    idu_rtu_rob_create_psrc2,
    idu_rtu_rob_create_dst,
    idu_rtu_rob_create_dst_vld,
    idu_rtu_rob_create_pdst,
    idu_rtu_rob_create_imm,
    idu_rtu_rob_create_imm_vld,
    idu_rtu_rob_create_type,
    idu_rtu_rob_create_pipe,
    idu_rtu_rob_create_ras,

    idu_rtu_rob_alu_issue_vld,
    idu_rtu_rob_alu_issue_iid,
    idu_rtu_rob_mxu_issue_vld,
    idu_rtu_rob_mxu_issue_iid,
    idu_rtu_rob_bju_issue_vld,
    idu_rtu_rob_bju_issue_iid,
    idu_rtu_rob_lsu_issue_vld,
    idu_rtu_rob_lsu_issue_iid,
    idu_rtu_rob_cp0_issue_vld,
    idu_rtu_rob_cp0_issue_iid,
    exu_rtu_rob_alu_complete_vld,
    exu_rtu_rob_alu_complete_iid,
    exu_rtu_rob_mxu_complete_vld,
    exu_rtu_rob_mxu_complete_iid,
    exu_rtu_rob_div_complete_vld,
    exu_rtu_rob_div_complete_iid,
    exu_rtu_rob_bju_complete_vld,
    exu_rtu_rob_bju_complete_iid,
    exu_rtu_rob_lsu_complete_vld,
    exu_rtu_rob_lsu_complete_iid,
    exu_rtu_rob_cp0_complete_vld,
    exu_rtu_rob_cp0_complete_iid,
    exu_rtu_rob_bju_pcjump_vld,
    exu_rtu_rob_bju_pcjump_iid,

    ebreak_gpr10,

    rtu_idu_rf_pcjump,
    rtu_global_flush,
    x_retire_vld,
    x_inst_retire_iid,

    iid_vld,
    iid
);
    // &Ports;
    input         clk;
    input         rst_clk;
    input         y_rtu_rob_stall_ctrl;
    input         idu_rtu_rob_iid_req_vld;
    input         idu_rtu_rob_create_vld;
    input  [6 :0] idu_rtu_rob_create_opcode;
    input  [2 :0] idu_rtu_rob_create_funct3;
    input  [63:0] idu_rtu_rob_create_pc;
    input  [4 :0] idu_rtu_rob_create_src1;
    input         idu_rtu_rob_create_src1_vld;
    input  [5 :0] idu_rtu_rob_create_psrc1;
    input  [4 :0] idu_rtu_rob_create_src2;
    input         idu_rtu_rob_create_src2_vld;
    input  [5 :0] idu_rtu_rob_create_psrc2;
    input  [4 :0] idu_rtu_rob_create_dst;
    input         idu_rtu_rob_create_dst_vld;
    input  [5 :0] idu_rtu_rob_create_pdst;
    input  [63:0] idu_rtu_rob_create_imm;
    input         idu_rtu_rob_create_imm_vld;
    input  [5 :0] idu_rtu_rob_create_type;
    input  [4 :0] idu_rtu_rob_create_pipe;
    input         idu_rtu_rob_create_ras;

    input         idu_rtu_rob_alu_issue_vld;
    input  [4 :0] idu_rtu_rob_alu_issue_iid;
    input         idu_rtu_rob_mxu_issue_vld;
    input  [4 :0] idu_rtu_rob_mxu_issue_iid;
    input         idu_rtu_rob_bju_issue_vld;
    input  [4 :0] idu_rtu_rob_bju_issue_iid;
    input         idu_rtu_rob_lsu_issue_vld;
    input  [4 :0] idu_rtu_rob_lsu_issue_iid;
    input         idu_rtu_rob_cp0_issue_vld;
    input  [4 :0] idu_rtu_rob_cp0_issue_iid;
    input         exu_rtu_rob_alu_complete_vld;
    input  [4 :0] exu_rtu_rob_alu_complete_iid;
    input         exu_rtu_rob_mxu_complete_vld;
    input  [4 :0] exu_rtu_rob_mxu_complete_iid;
    input         exu_rtu_rob_div_complete_vld;
    input  [4 :0] exu_rtu_rob_div_complete_iid;
    input         exu_rtu_rob_bju_complete_vld;
    input  [4 :0] exu_rtu_rob_bju_complete_iid;
    input         exu_rtu_rob_lsu_complete_vld;
    input  [4 :0] exu_rtu_rob_lsu_complete_iid;
    input         exu_rtu_rob_cp0_complete_vld;
    input  [4 :0] exu_rtu_rob_cp0_complete_iid;
    input         exu_rtu_rob_bju_pcjump_vld;
    input  [4 :0] exu_rtu_rob_bju_pcjump_iid;

    input  [63:0] ebreak_gpr10;

    output        rtu_idu_rf_pcjump;
    output        rtu_global_flush;
    output        x_retire_vld;
    output [4 :0] x_inst_retire_iid;

    output        iid_vld;
    output [4 :0] iid;

    // &Regs;
    reg [4 :0] head_iid_ptr;
    reg [4 :0] tail_iid_ptr;
    reg [4 :0] num;

    // &Wires;
    wire        clk;
    wire        rst_clk;
    wire        y_rtu_rob_stall_ctrl;
    wire        idu_rtu_rob_iid_req_vld;
    wire        idu_rtu_rob_create_vld;
    wire [6 :0] idu_rtu_rob_create_opcode;
    wire [2 :0] idu_rtu_rob_create_funct3;
    wire [63:0] idu_rtu_rob_create_pc;
    wire [4 :0] idu_rtu_rob_create_src1;
    wire        idu_rtu_rob_create_src1_vld;
    wire [5 :0] idu_rtu_rob_create_psrc1;
    wire [4 :0] idu_rtu_rob_create_src2;
    wire        idu_rtu_rob_create_src2_vld;
    wire [5 :0] idu_rtu_rob_create_psrc2;
    wire [4 :0] idu_rtu_rob_create_dst;
    wire        idu_rtu_rob_create_dst_vld;
    wire [5 :0] idu_rtu_rob_create_pdst;
    wire [63:0] idu_rtu_rob_create_imm;
    wire        idu_rtu_rob_create_imm_vld;
    wire [5 :0] idu_rtu_rob_create_type;
    wire [4 :0] idu_rtu_rob_create_pipe;
    wire        idu_rtu_rob_create_ras;

    wire        idu_rtu_rob_alu_issue_vld;
    wire [4 :0] idu_rtu_rob_alu_issue_iid;
    wire        idu_rtu_rob_mxu_issue_vld;
    wire [4 :0] idu_rtu_rob_mxu_issue_iid;
    wire        idu_rtu_rob_bju_issue_vld;
    wire [4 :0] idu_rtu_rob_bju_issue_iid;
    wire        idu_rtu_rob_lsu_issue_vld;
    wire [4 :0] idu_rtu_rob_lsu_issue_iid;
    wire        idu_rtu_rob_cp0_issue_vld;
    wire [4 :0] idu_rtu_rob_cp0_issue_iid;
    wire        exu_rtu_rob_alu_complete_vld;
    wire [4 :0] exu_rtu_rob_alu_complete_iid;
    wire        exu_rtu_rob_mxu_complete_vld;
    wire [4 :0] exu_rtu_rob_mxu_complete_iid;
    wire        exu_rtu_rob_div_complete_vld;
    wire [4 :0] exu_rtu_rob_div_complete_iid;
    wire        exu_rtu_rob_bju_complete_vld;
    wire [4 :0] exu_rtu_rob_bju_complete_iid;
    wire        exu_rtu_rob_lsu_complete_vld;
    wire [4 :0] exu_rtu_rob_lsu_complete_iid;
    wire        exu_rtu_rob_cp0_complete_vld;
    wire [4 :0] exu_rtu_rob_cp0_complete_iid;
    wire        exu_rtu_rob_bju_pcjump_vld;
    wire [4 :0] exu_rtu_rob_bju_pcjump_iid;

    wire [63:0] ebreak_gpr10;

    wire        rtu_idu_rf_pcjump;
    wire        rtu_global_flush;
    wire        x_retire_vld;
    wire [4 :0] x_inst_retire_iid;
    wire        iid_invalid;
    wire        iid_vld;
    wire [4 :0] iid;
    wire        rob_full_stats;
    wire        rob_empty_stats;
    wire        rob_create_vld;
    wire        rob_retire_vld;
    wire [15:0] create_vld;
    wire [15:0] head_iid_ptr_cur_vld;
    wire [15:0] retire_vld;
    wire [15:0] jump_vld;
    wire [15:0] flush_vld;
    wire [15:0] issue_vld;
    wire [15:0] complete_vld;
    wire [15:0] bju_vld;

    wire [190:0] iid0_message;
    wire [190:0] iid1_message;
    wire [190:0] iid2_message;
    wire [190:0] iid3_message;
    wire [190:0] iid4_message;
    wire [190:0] iid5_message;
    wire [190:0] iid6_message;
    wire [190:0] iid7_message;
    wire [190:0] iid8_message;
    wire [190:0] iid9_message;
    wire [190:0] iid10_message;
    wire [190:0] iid11_message;
    wire [190:0] iid12_message;
    wire [190:0] iid13_message;
    wire [190:0] iid14_message;
    wire [190:0] iid15_message;

    rtu_rob_entry rtu_rob_iid0_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[0]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[0]               ),
        .complete_vld           (complete_vld[0]            ),
        .bju_vld                (bju_vld[0]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[0]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[0]              ),
        .jump_vld               (jump_vld[0]                ),
        .flush_vld              (flush_vld[0]               ),
        .inst_message           (iid0_message               )
    );

    rtu_rob_entry rtu_rob_iid1_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[1]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[1]               ),
        .complete_vld           (complete_vld[1]            ),
        .bju_vld                (bju_vld[1]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[1]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[1]              ),
        .jump_vld               (jump_vld[1]                ),
        .flush_vld              (flush_vld[1]               ),
        .inst_message           (iid1_message               )
    );

    rtu_rob_entry rtu_rob_iid2_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[2]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[2]               ),
        .complete_vld           (complete_vld[2]            ),
        .bju_vld                (bju_vld[2]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[2]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[2]              ),
        .jump_vld               (jump_vld[2]                ),
        .flush_vld              (flush_vld[2]               ),
        .inst_message           (iid2_message               )
    );

    rtu_rob_entry rtu_rob_iid3_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[3]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[3]               ),
        .complete_vld           (complete_vld[3]            ),
        .bju_vld                (bju_vld[3]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[3]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[3]              ),
        .jump_vld               (jump_vld[3]                ),
        .flush_vld              (flush_vld[3]               ),
        .inst_message           (iid3_message               )
    );

    rtu_rob_entry rtu_rob_iid4_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[4]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[4]               ),
        .complete_vld           (complete_vld[4]            ),
        .bju_vld                (bju_vld[4]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[4]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[4]              ),
        .jump_vld               (jump_vld[4]                ),
        .flush_vld              (flush_vld[4]               ),
        .inst_message           (iid4_message               )
    );

    rtu_rob_entry rtu_rob_iid5_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[5]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[5]               ),
        .complete_vld           (complete_vld[5]            ),
        .bju_vld                (bju_vld[5]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[5]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[5]              ),
        .jump_vld               (jump_vld[5]                ),
        .flush_vld              (flush_vld[5]               ),
        .inst_message           (iid5_message               )
    );

    rtu_rob_entry rtu_rob_iid6_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[6]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[6]               ),
        .complete_vld           (complete_vld[6]            ),
        .bju_vld                (bju_vld[6]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[6]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[6]              ),
        .jump_vld               (jump_vld[6]                ),
        .flush_vld              (flush_vld[6]               ),
        .inst_message           (iid6_message               )
    );

    rtu_rob_entry rtu_rob_iid7_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[7]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[7]               ),
        .complete_vld           (complete_vld[7]            ),
        .bju_vld                (bju_vld[7]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[7]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[7]              ),
        .jump_vld               (jump_vld[7]                ),
        .flush_vld              (flush_vld[7]               ),
        .inst_message           (iid7_message               )
    );

    rtu_rob_entry rtu_rob_iid8_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[8]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[8]               ),
        .complete_vld           (complete_vld[8]            ),
        .bju_vld                (bju_vld[8]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[8]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[8]              ),
        .jump_vld               (jump_vld[8]                ),
        .flush_vld              (flush_vld[8]               ),
        .inst_message           (iid8_message               )
    );

    rtu_rob_entry rtu_rob_iid9_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[9]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[9]               ),
        .complete_vld           (complete_vld[9]            ),
        .bju_vld                (bju_vld[9]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[9]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[9]              ),
        .jump_vld               (jump_vld[9]                ),
        .flush_vld              (flush_vld[9]               ),
        .inst_message           (iid9_message               )
    );

    rtu_rob_entry rtu_rob_iid10_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[10]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[10]               ),
        .complete_vld           (complete_vld[10]            ),
        .bju_vld                (bju_vld[10]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[10]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[10]              ),
        .jump_vld               (jump_vld[10]                ),
        .flush_vld              (flush_vld[10]               ),
        .inst_message           (iid10_message               )
    );

    rtu_rob_entry rtu_rob_iid11_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[11]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[11]               ),
        .complete_vld           (complete_vld[11]            ),
        .bju_vld                (bju_vld[11]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[11]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[11]              ),
        .jump_vld               (jump_vld[11]                ),
        .flush_vld              (flush_vld[11]               ),
        .inst_message           (iid11_message               )
    );

    rtu_rob_entry rtu_rob_iid12_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[12]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[12]               ),
        .complete_vld           (complete_vld[12]            ),
        .bju_vld                (bju_vld[12]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[12]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[12]              ),
        .jump_vld               (jump_vld[12]                ),
        .flush_vld              (flush_vld[12]               ),
        .inst_message           (iid12_message               )
    );

    rtu_rob_entry rtu_rob_iid13_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[13]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[13]               ),
        .complete_vld           (complete_vld[13]            ),
        .bju_vld                (bju_vld[13]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[13]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[13]              ),
        .jump_vld               (jump_vld[13]                ),
        .flush_vld              (flush_vld[13]               ),
        .inst_message           (iid13_message               )
    );

    rtu_rob_entry rtu_rob_iid14_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[14]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[14]               ),
        .complete_vld           (complete_vld[14]            ),
        .bju_vld                (bju_vld[14]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[14]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[14]              ),
        .jump_vld               (jump_vld[14]                ),
        .flush_vld              (flush_vld[14]               ),
        .inst_message           (iid14_message               )
    );

    rtu_rob_entry rtu_rob_iid15_entry(
        .clk                    (clk                            ),
        .rst_clk                (rst_clk                        ),
        .create_vld             (create_vld[15]              ),
        .create_opcode          (idu_rtu_rob_create_opcode      ),
        .create_funct3          (idu_rtu_rob_create_funct3      ),
        .create_pc              (idu_rtu_rob_create_pc          ),
        .create_src1            (idu_rtu_rob_create_src1        ),
        .create_src1_vld        (idu_rtu_rob_create_src1_vld    ),
        .create_psrc1           (idu_rtu_rob_create_psrc1       ),
        .create_src2            (idu_rtu_rob_create_src2        ),
        .create_src2_vld        (idu_rtu_rob_create_src2_vld    ),
        .create_psrc2           (idu_rtu_rob_create_psrc2       ),
        .create_dst             (idu_rtu_rob_create_dst         ),
        .create_dst_vld         (idu_rtu_rob_create_dst_vld     ),
        .create_pdst            (idu_rtu_rob_create_pdst        ),
        .create_imm             (idu_rtu_rob_create_imm         ),
        .create_imm_vld         (idu_rtu_rob_create_imm_vld     ),
        .create_type            (idu_rtu_rob_create_type        ),
        .create_pipe            (idu_rtu_rob_create_pipe        ),
        .create_ras             (idu_rtu_rob_create_ras         ),
        .issue_vld              (issue_vld[15]               ),
        .complete_vld           (complete_vld[15]            ),
        .bju_vld                (bju_vld[15]                 ),
        .rtu_global_flush       (rtu_global_flush               ),
        .head_iid_ptr_cur_vld   (head_iid_ptr_cur_vld[15]    ),
        .ebreak_gpr10           (ebreak_gpr10                   ),
        .retire_vld             (retire_vld[15]              ),
        .jump_vld               (jump_vld[15]                ),
        .flush_vld              (flush_vld[15]               ),
        .inst_message           (iid15_message               )
    );

    // issue sign
    for (genvar i = 0; i < 16; i++)
    begin: issue_sign
        assign issue_vld[i] = (idu_rtu_rob_alu_issue_vld & (idu_rtu_rob_alu_issue_iid[3:0] == i))
                            | (idu_rtu_rob_mxu_issue_vld & (idu_rtu_rob_mxu_issue_iid[3:0] == i))
                            | (idu_rtu_rob_bju_issue_vld & (idu_rtu_rob_bju_issue_iid[3:0] == i))
                            | (idu_rtu_rob_lsu_issue_vld & (idu_rtu_rob_lsu_issue_iid[3:0] == i))
                            | (idu_rtu_rob_cp0_issue_vld & (idu_rtu_rob_cp0_issue_iid[3:0] == i));
    end

    // complete sign
    for (genvar i = 0; i < 16; i++)
    begin: complete_sign
        assign complete_vld[i] = (exu_rtu_rob_alu_complete_vld & (exu_rtu_rob_alu_complete_iid[3:0] == i))
                               | (exu_rtu_rob_mxu_complete_vld & (exu_rtu_rob_mxu_complete_iid[3:0] == i))
                               | (exu_rtu_rob_div_complete_vld & (exu_rtu_rob_div_complete_iid[3:0] == i))
                               | (exu_rtu_rob_bju_complete_vld & (exu_rtu_rob_bju_complete_iid[3:0] == i))
                               | (exu_rtu_rob_lsu_complete_vld & (exu_rtu_rob_lsu_complete_iid[3:0] == i))
                               | (exu_rtu_rob_cp0_complete_vld & (exu_rtu_rob_cp0_complete_iid[3:0] == i));
    end

    // bju_vld_sign
    for (genvar i = 0; i < 16; i++)
    begin: bju_sign
        assign bju_vld[i] = exu_rtu_rob_bju_pcjump_vld & (exu_rtu_rob_bju_pcjump_iid[3:0] == i);
    end

    // iid req
    assign rob_full_stats = (num == 16);
    assign iid_invalid    = idu_rtu_rob_iid_req_vld || !iid_vld;
    assign iid_vld        = !rob_full_stats;

    // iid create
    assign rob_create_vld = idu_rtu_rob_create_vld & !rob_full_stats & ~y_rtu_rob_stall_ctrl;
    assign iid            = tail_iid_ptr;
    for (genvar i = 0; i < 16; i++)
    begin: create_vld_sign
        assign create_vld[i] = (tail_iid_ptr[3:0] == i) & rob_create_vld;
    end

    always @(posedge clk or negedge rst_clk)
    begin
        if (!rst_clk)
            tail_iid_ptr <= 5'b0;
        else if (rtu_global_flush)
            tail_iid_ptr <= 5'b0;
        else if (rob_create_vld)
            tail_iid_ptr <= tail_iid_ptr + 1;
        else
            tail_iid_ptr <= tail_iid_ptr;
    end

    // iid pop
    assign rob_empty_stats   = (num == 0);
    assign x_retire_vld      = |retire_vld[15:0];
    assign x_inst_retire_iid = head_iid_ptr;
    assign rob_retire_vld = x_retire_vld & !rob_empty_stats;
    for (genvar i = 0; i < 16; i++)
    begin: head_iid_ptr_cur_vld_sign
        assign head_iid_ptr_cur_vld[i] = (head_iid_ptr[3:0] == i);
    end

    always @(posedge clk or negedge rst_clk)
    begin
        if (!rst_clk)
            head_iid_ptr <= 5'b0;
        else if (rtu_global_flush)
            head_iid_ptr <= 5'b0;
        else if (rob_retire_vld)
            head_iid_ptr <= head_iid_ptr + 1;
        else
            head_iid_ptr <= head_iid_ptr;
    end

    // num
    always @(posedge clk or negedge rst_clk)
    begin
        if (!rst_clk)
            num <= 0;
        else if (rtu_global_flush)
            num <= 0;
        else if (rob_create_vld && rob_retire_vld)
            num <= num;
        else if (rob_create_vld)
            num <= num + 1;
        else if (rob_retire_vld)
            num <= num - 1;
        else
            num <= num;
    end

    // jump and flush
    assign rtu_idu_rf_pcjump = |jump_vld[15:0];
    assign rtu_global_flush = |flush_vld[15:0];

    // DEBUG for Prove Out-of-Order
    `ifdef DEBUG_RTU_ROB_PRINT
        always @(negedge clk)
        begin: message_print
            $display("RTU_ROB: iid = %d, vld = %b, num = %d", iid, iid_vld, num);
            $display("|                                                 |    jump   |           src1          |           src2          |          dst         |            imm             |  type  |            pipe             |       stats        |");
            $display("| iid | vld | opcode  | funct3 |        pc        | bju | ras | src1_vld | src1 | psrc1 | src2_vld | src2 | psrc2 | dst_vld | dst | pdst | imm_vld |       imm        | RISBUJ | ALU | MXU | BJU | LSU | CP0 | issue? | complete? |");
            $display("| 0   | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid0_message[190],     iid0_message[189:183], iid0_message[182:180], iid0_message[179:116],
                    iid0_message[115],     iid0_message[114],     iid0_message[113],     iid0_message[112:108],
                    iid0_message[107:102], iid0_message[101],     iid0_message[100:96],  iid0_message[95:90],
                    iid0_message[89],      iid0_message[88:84],   iid0_message[83:78],   iid0_message[77],
                    iid0_message[76:13],   iid0_message[12:7],    iid0_message[6],       iid0_message[5],
                    iid0_message[4],       iid0_message[3],       iid0_message[2],       iid0_message[1],       iid0_message[0]);
            $display("| 1   | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid1_message[190],     iid1_message[189:183], iid1_message[182:180], iid1_message[179:116],
                    iid1_message[115],     iid1_message[114],     iid1_message[113],     iid1_message[112:108],
                    iid1_message[107:102], iid1_message[101],     iid1_message[100:96],  iid1_message[95:90],
                    iid1_message[89],      iid1_message[88:84],   iid1_message[83:78],   iid1_message[77],
                    iid1_message[76:13],   iid1_message[12:7],    iid1_message[6],       iid1_message[5],
                    iid1_message[4],       iid1_message[3],       iid1_message[2],       iid1_message[1],       iid1_message[0]);
            $display("| 2   | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid2_message[190],     iid2_message[189:183], iid2_message[182:180], iid2_message[179:116],
                    iid2_message[115],     iid2_message[114],     iid2_message[113],     iid2_message[112:108],
                    iid2_message[107:102], iid2_message[101],     iid2_message[100:96],  iid2_message[95:90],
                    iid2_message[89],      iid2_message[88:84],   iid2_message[83:78],   iid2_message[77],
                    iid2_message[76:13],   iid2_message[12:7],    iid2_message[6],       iid2_message[5],
                    iid2_message[4],       iid2_message[3],       iid2_message[2],       iid2_message[1],       iid2_message[0]);
            $display("| 3   | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid3_message[190],     iid3_message[189:183], iid3_message[182:180], iid3_message[179:116],
                    iid3_message[115],     iid3_message[114],     iid3_message[113],     iid3_message[112:108],
                    iid3_message[107:102], iid3_message[101],     iid3_message[100:96],  iid3_message[95:90],
                    iid3_message[89],      iid3_message[88:84],   iid3_message[83:78],   iid3_message[77],
                    iid3_message[76:13],   iid3_message[12:7],    iid3_message[6],       iid3_message[5],
                    iid3_message[4],       iid3_message[3],       iid3_message[2],       iid3_message[1],       iid3_message[0]);
            $display("| 4   | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid4_message[190],     iid4_message[189:183], iid4_message[182:180], iid4_message[179:116],
                    iid4_message[115],     iid4_message[114],     iid4_message[113],     iid4_message[112:108],
                    iid4_message[107:102], iid4_message[101],     iid4_message[100:96],  iid4_message[95:90],
                    iid4_message[89],      iid4_message[88:84],   iid4_message[83:78],   iid4_message[77],
                    iid4_message[76:13],   iid4_message[12:7],    iid4_message[6],       iid4_message[5],
                    iid4_message[4],       iid4_message[3],       iid4_message[2],       iid4_message[1],       iid4_message[0]);
            $display("| 5   | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid5_message[190],     iid5_message[189:183], iid5_message[182:180], iid5_message[179:116],
                    iid5_message[115],     iid5_message[114],     iid5_message[113],     iid5_message[112:108],
                    iid5_message[107:102], iid5_message[101],     iid5_message[100:96],  iid5_message[95:90],
                    iid5_message[89],      iid5_message[88:84],   iid5_message[83:78],   iid5_message[77],
                    iid5_message[76:13],   iid5_message[12:7],    iid5_message[6],       iid5_message[5],
                    iid5_message[4],       iid5_message[3],       iid5_message[2],       iid5_message[1],       iid5_message[0]);
            $display("| 6   | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid6_message[190],     iid6_message[189:183], iid6_message[182:180], iid6_message[179:116],
                    iid6_message[115],     iid6_message[114],     iid6_message[113],     iid6_message[112:108],
                    iid6_message[107:102], iid6_message[101],     iid6_message[100:96],  iid6_message[95:90],
                    iid6_message[89],      iid6_message[88:84],   iid6_message[83:78],   iid6_message[77],
                    iid6_message[76:13],   iid6_message[12:7],    iid6_message[6],       iid6_message[5],
                    iid6_message[4],       iid6_message[3],       iid6_message[2],       iid6_message[1],       iid6_message[0]);
            $display("| 7   | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid7_message[190],     iid7_message[189:183], iid7_message[182:180], iid7_message[179:116],
                    iid7_message[115],     iid7_message[114],     iid7_message[113],     iid7_message[112:108],
                    iid7_message[107:102], iid7_message[101],     iid7_message[100:96],  iid7_message[95:90],
                    iid7_message[89],      iid7_message[88:84],   iid7_message[83:78],   iid7_message[77],
                    iid7_message[76:13],   iid7_message[12:7],    iid7_message[6],       iid7_message[5],
                    iid7_message[4],       iid7_message[3],       iid7_message[2],       iid7_message[1],       iid7_message[0]);
            $display("| 8   | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid8_message[190],     iid8_message[189:183], iid8_message[182:180], iid8_message[179:116],
                    iid8_message[115],     iid8_message[114],     iid8_message[113],     iid8_message[112:108],
                    iid8_message[107:102], iid8_message[101],     iid8_message[100:96],  iid8_message[95:90],
                    iid8_message[89],      iid8_message[88:84],   iid8_message[83:78],   iid8_message[77],
                    iid8_message[76:13],   iid8_message[12:7],    iid8_message[6],       iid8_message[5],
                    iid8_message[4],       iid8_message[3],       iid8_message[2],       iid8_message[1],       iid8_message[0]);
            $display("| 9   | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid9_message[190],     iid9_message[189:183], iid9_message[182:180], iid9_message[179:116],
                    iid9_message[115],     iid9_message[114],     iid9_message[113],     iid9_message[112:108],
                    iid9_message[107:102], iid9_message[101],     iid9_message[100:96],  iid9_message[95:90],
                    iid9_message[89],      iid9_message[88:84],   iid9_message[83:78],   iid9_message[77],
                    iid9_message[76:13],   iid9_message[12:7],    iid9_message[6],       iid9_message[5],
                    iid9_message[4],       iid9_message[3],       iid9_message[2],       iid9_message[1],       iid9_message[0]);
            $display("| 10  | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid10_message[190],     iid10_message[189:183], iid10_message[182:180], iid10_message[179:116],
                    iid10_message[115],     iid10_message[114],     iid10_message[113],     iid10_message[112:108],
                    iid10_message[107:102], iid10_message[101],     iid10_message[100:96],  iid10_message[95:90],
                    iid10_message[89],      iid10_message[88:84],   iid10_message[83:78],   iid10_message[77],
                    iid10_message[76:13],   iid10_message[12:7],    iid10_message[6],       iid10_message[5],
                    iid10_message[4],       iid10_message[3],       iid10_message[2],       iid10_message[1],       iid10_message[0]);
            $display("| 11  | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid11_message[190],     iid11_message[189:183], iid11_message[182:180], iid11_message[179:116],
                    iid11_message[115],     iid11_message[114],     iid11_message[113],     iid11_message[112:108],
                    iid11_message[107:102], iid11_message[101],     iid11_message[100:96],  iid11_message[95:90],
                    iid11_message[89],      iid11_message[88:84],   iid11_message[83:78],   iid11_message[77],
                    iid11_message[76:13],   iid11_message[12:7],    iid11_message[6],       iid11_message[5],
                    iid11_message[4],       iid11_message[3],       iid11_message[2],       iid11_message[1],       iid11_message[0]);
            $display("| 12  | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid12_message[190],     iid12_message[189:183], iid12_message[182:180], iid12_message[179:116],
                    iid12_message[115],     iid12_message[114],     iid12_message[113],     iid12_message[112:108],
                    iid12_message[107:102], iid12_message[101],     iid12_message[100:96],  iid12_message[95:90],
                    iid12_message[89],      iid12_message[88:84],   iid12_message[83:78],   iid12_message[77],
                    iid12_message[76:13],   iid12_message[12:7],    iid12_message[6],       iid12_message[5],
                    iid12_message[4],       iid12_message[3],       iid12_message[2],       iid12_message[1],       iid12_message[0]);
            $display("| 13  | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid13_message[190],     iid13_message[189:183], iid13_message[182:180], iid13_message[179:116],
                    iid13_message[115],     iid13_message[114],     iid13_message[113],     iid13_message[112:108],
                    iid13_message[107:102], iid13_message[101],     iid13_message[100:96],  iid13_message[95:90],
                    iid13_message[89],      iid13_message[88:84],   iid13_message[83:78],   iid13_message[77],
                    iid13_message[76:13],   iid13_message[12:7],    iid13_message[6],       iid13_message[5],
                    iid13_message[4],       iid13_message[3],       iid13_message[2],       iid13_message[1],       iid13_message[0]);
            $display("| 14  | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid14_message[190],     iid14_message[189:183], iid14_message[182:180], iid14_message[179:116],
                    iid14_message[115],     iid14_message[114],     iid14_message[113],     iid14_message[112:108],
                    iid14_message[107:102], iid14_message[101],     iid14_message[100:96],  iid14_message[95:90],
                    iid14_message[89],      iid14_message[88:84],   iid14_message[83:78],   iid14_message[77],
                    iid14_message[76:13],   iid14_message[12:7],    iid14_message[6],       iid14_message[5],
                    iid14_message[4],       iid14_message[3],       iid14_message[2],       iid14_message[1],       iid14_message[0]);
            $display("| 15  | %b   | %b | %b    | %x | %b   | %b   | %b        | x%02d  | p%02d   | %b        | x%02d  | p%02d   | %b       | x%02d | p%02d  | %b       | %x | %b | %b   | %b   | %b   | %b   | %b   | %b      | %b         |",
                    iid15_message[190],     iid15_message[189:183], iid15_message[182:180], iid15_message[179:116],
                    iid15_message[115],     iid15_message[114],     iid15_message[113],     iid15_message[112:108],
                    iid15_message[107:102], iid15_message[101],     iid15_message[100:96],  iid15_message[95:90],
                    iid15_message[89],      iid15_message[88:84],   iid15_message[83:78],   iid15_message[77],
                    iid15_message[76:13],   iid15_message[12:7],    iid15_message[6],       iid15_message[5],
                    iid15_message[4],       iid15_message[3],       iid15_message[2],       iid15_message[1],       iid15_message[0]);
        end
    `endif

endmodule
