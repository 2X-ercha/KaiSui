module rtu_pst_preg (
    clk,
    rst_clk,
    rtu_global_flush,
    idu_rtu_pst_pdst_req_vld,
    idu_rtu_pst_create_vld,
    idu_rtu_pst_create_preg_index,
    idu_rtu_pst_create_iid,
    idu_rtu_pst_create_gpr_index,
    idu_rtu_pst_create_gpr_pre_preg_index,
    x_inst_retire_iid,
    x_retire_vld,
    idu_rtu_pst_wb_vld,
    alloc_preg_vld,
    alloc_preg,
    rtu_idu_ir_recover_table
);
    // &Ports;
    input         clk;
    input         rst_clk;
    input         rtu_global_flush;
    input         idu_rtu_pst_pdst_req_vld;
    input         idu_rtu_pst_create_vld;
    input  [5 :0] idu_rtu_pst_create_preg_index;
    input  [3 :0] idu_rtu_pst_create_iid;
    input  [4 :0] idu_rtu_pst_create_gpr_index;
    input  [5 :0] idu_rtu_pst_create_gpr_pre_preg_index;
    input  [3 :0] x_inst_retire_iid;
    input         x_retire_vld;
    input  [63:0] idu_rtu_pst_wb_vld;
    output        alloc_preg_vld;
    output [5 :0] alloc_preg;
    output [191:0] rtu_idu_ir_recover_table;

    // &Regs;
    reg        alloc_preg_vld;
    reg [5 :0] alloc_preg;

    // &Wires;
    wire        clk;
    wire        rst_clk;
    wire        rtu_global_flush;
    wire        idu_rtu_pst_pdst_req_vld;
    wire        idu_rtu_pst_create_vld;
    wire [3 :0] idu_rtu_pst_create_iid;
    wire [4 :0] idu_rtu_pst_create_gpr_index;
    wire [5 :0] idu_rtu_pst_create_gpr_pre_preg_index;
    wire [3 :0] x_inst_retire_iid;
    wire        x_retire_vld;
    wire [63:0] idu_rtu_pst_wb_vld;
    wire [191:0] rtu_idu_ir_recover_table;

    wire [63:0] preg_dealloc;
    wire [63:0] preg_pre_alloc_priority;
    wire [63:0] preg_pre_alloc_vld;
    wire [5 :0] pre_alloc_preg;
    wire [63:0] preg_alloc_vld;
    wire        alloc_preg_invalid;
    wire        pre_alloc_vld;
    wire [63:0] preg_release_vld;
    wire [63:0] preg0_release_expand;
    wire [63:0] preg1_release_expand;
    wire [63:0] preg2_release_expand;
    wire [63:0] preg3_release_expand;
    wire [63:0] preg4_release_expand;
    wire [63:0] preg5_release_expand;
    wire [63:0] preg6_release_expand;
    wire [63:0] preg7_release_expand;
    wire [63:0] preg8_release_expand;
    wire [63:0] preg9_release_expand;
    wire [63:0] preg10_release_expand;
    wire [63:0] preg11_release_expand;
    wire [63:0] preg12_release_expand;
    wire [63:0] preg13_release_expand;
    wire [63:0] preg14_release_expand;
    wire [63:0] preg15_release_expand;
    wire [63:0] preg16_release_expand;
    wire [63:0] preg17_release_expand;
    wire [63:0] preg18_release_expand;
    wire [63:0] preg19_release_expand;
    wire [63:0] preg20_release_expand;
    wire [63:0] preg21_release_expand;
    wire [63:0] preg22_release_expand;
    wire [63:0] preg23_release_expand;
    wire [63:0] preg24_release_expand;
    wire [63:0] preg25_release_expand;
    wire [63:0] preg26_release_expand;
    wire [63:0] preg27_release_expand;
    wire [63:0] preg28_release_expand;
    wire [63:0] preg29_release_expand;
    wire [63:0] preg30_release_expand;
    wire [63:0] preg31_release_expand;
    wire [63:0] preg32_release_expand;
    wire [63:0] preg33_release_expand;
    wire [63:0] preg34_release_expand;
    wire [63:0] preg35_release_expand;
    wire [63:0] preg36_release_expand;
    wire [63:0] preg37_release_expand;
    wire [63:0] preg38_release_expand;
    wire [63:0] preg39_release_expand;
    wire [63:0] preg40_release_expand;
    wire [63:0] preg41_release_expand;
    wire [63:0] preg42_release_expand;
    wire [63:0] preg43_release_expand;
    wire [63:0] preg44_release_expand;
    wire [63:0] preg45_release_expand;
    wire [63:0] preg46_release_expand;
    wire [63:0] preg47_release_expand;
    wire [63:0] preg48_release_expand;
    wire [63:0] preg49_release_expand;
    wire [63:0] preg50_release_expand;
    wire [63:0] preg51_release_expand;
    wire [63:0] preg52_release_expand;
    wire [63:0] preg53_release_expand;
    wire [63:0] preg54_release_expand;
    wire [63:0] preg55_release_expand;
    wire [63:0] preg56_release_expand;
    wire [63:0] preg57_release_expand;
    wire [63:0] preg58_release_expand;
    wire [63:0] preg59_release_expand;
    wire [63:0] preg60_release_expand;
    wire [63:0] preg61_release_expand;
    wire [63:0] preg62_release_expand;
    wire [63:0] preg63_release_expand;
    wire [63:0] preg_reset_mapped;
    // wire [4 :0] preg0_reset_gpr_mapped;
    wire [4 :0] preg1_reset_gpr_mapped;
    wire [4 :0] preg2_reset_gpr_mapped;
    wire [4 :0] preg3_reset_gpr_mapped;
    wire [4 :0] preg4_reset_gpr_mapped;
    wire [4 :0] preg5_reset_gpr_mapped;
    wire [4 :0] preg6_reset_gpr_mapped;
    wire [4 :0] preg7_reset_gpr_mapped;
    wire [4 :0] preg8_reset_gpr_mapped;
    wire [4 :0] preg9_reset_gpr_mapped;
    wire [4 :0] preg10_reset_gpr_mapped;
    wire [4 :0] preg11_reset_gpr_mapped;
    wire [4 :0] preg12_reset_gpr_mapped;
    wire [4 :0] preg13_reset_gpr_mapped;
    wire [4 :0] preg14_reset_gpr_mapped;
    wire [4 :0] preg15_reset_gpr_mapped;
    wire [4 :0] preg16_reset_gpr_mapped;
    wire [4 :0] preg17_reset_gpr_mapped;
    wire [4 :0] preg18_reset_gpr_mapped;
    wire [4 :0] preg19_reset_gpr_mapped;
    wire [4 :0] preg20_reset_gpr_mapped;
    wire [4 :0] preg21_reset_gpr_mapped;
    wire [4 :0] preg22_reset_gpr_mapped;
    wire [4 :0] preg23_reset_gpr_mapped;
    wire [4 :0] preg24_reset_gpr_mapped;
    wire [4 :0] preg25_reset_gpr_mapped;
    wire [4 :0] preg26_reset_gpr_mapped;
    wire [4 :0] preg27_reset_gpr_mapped;
    wire [4 :0] preg28_reset_gpr_mapped;
    wire [4 :0] preg29_reset_gpr_mapped;
    wire [4 :0] preg30_reset_gpr_mapped;
    wire [4 :0] preg31_reset_gpr_mapped;
    wire [4 :0] preg32_reset_gpr_mapped;
    wire [4 :0] preg33_reset_gpr_mapped;
    wire [4 :0] preg34_reset_gpr_mapped;
    wire [4 :0] preg35_reset_gpr_mapped;
    wire [4 :0] preg36_reset_gpr_mapped;
    wire [4 :0] preg37_reset_gpr_mapped;
    wire [4 :0] preg38_reset_gpr_mapped;
    wire [4 :0] preg39_reset_gpr_mapped;
    wire [4 :0] preg40_reset_gpr_mapped;
    wire [4 :0] preg41_reset_gpr_mapped;
    wire [4 :0] preg42_reset_gpr_mapped;
    wire [4 :0] preg43_reset_gpr_mapped;
    wire [4 :0] preg44_reset_gpr_mapped;
    wire [4 :0] preg45_reset_gpr_mapped;
    wire [4 :0] preg46_reset_gpr_mapped;
    wire [4 :0] preg47_reset_gpr_mapped;
    wire [4 :0] preg48_reset_gpr_mapped;
    wire [4 :0] preg49_reset_gpr_mapped;
    wire [4 :0] preg50_reset_gpr_mapped;
    wire [4 :0] preg51_reset_gpr_mapped;
    wire [4 :0] preg52_reset_gpr_mapped;
    wire [4 :0] preg53_reset_gpr_mapped;
    wire [4 :0] preg54_reset_gpr_mapped;
    wire [4 :0] preg55_reset_gpr_mapped;
    wire [4 :0] preg56_reset_gpr_mapped;
    wire [4 :0] preg57_reset_gpr_mapped;
    wire [4 :0] preg58_reset_gpr_mapped;
    wire [4 :0] preg59_reset_gpr_mapped;
    wire [4 :0] preg60_reset_gpr_mapped;
    wire [4 :0] preg61_reset_gpr_mapped;
    wire [4 :0] preg62_reset_gpr_mapped;
    wire [4 :0] preg63_reset_gpr_mapped;
    wire [31:0] preg0_recover_table_to_gpr;
    wire [31:0] preg1_recover_table_to_gpr;
    wire [31:0] preg2_recover_table_to_gpr;
    wire [31:0] preg3_recover_table_to_gpr;
    wire [31:0] preg4_recover_table_to_gpr;
    wire [31:0] preg5_recover_table_to_gpr;
    wire [31:0] preg6_recover_table_to_gpr;
    wire [31:0] preg7_recover_table_to_gpr;
    wire [31:0] preg8_recover_table_to_gpr;
    wire [31:0] preg9_recover_table_to_gpr;
    wire [31:0] preg10_recover_table_to_gpr;
    wire [31:0] preg11_recover_table_to_gpr;
    wire [31:0] preg12_recover_table_to_gpr;
    wire [31:0] preg13_recover_table_to_gpr;
    wire [31:0] preg14_recover_table_to_gpr;
    wire [31:0] preg15_recover_table_to_gpr;
    wire [31:0] preg16_recover_table_to_gpr;
    wire [31:0] preg17_recover_table_to_gpr;
    wire [31:0] preg18_recover_table_to_gpr;
    wire [31:0] preg19_recover_table_to_gpr;
    wire [31:0] preg20_recover_table_to_gpr;
    wire [31:0] preg21_recover_table_to_gpr;
    wire [31:0] preg22_recover_table_to_gpr;
    wire [31:0] preg23_recover_table_to_gpr;
    wire [31:0] preg24_recover_table_to_gpr;
    wire [31:0] preg25_recover_table_to_gpr;
    wire [31:0] preg26_recover_table_to_gpr;
    wire [31:0] preg27_recover_table_to_gpr;
    wire [31:0] preg28_recover_table_to_gpr;
    wire [31:0] preg29_recover_table_to_gpr;
    wire [31:0] preg30_recover_table_to_gpr;
    wire [31:0] preg31_recover_table_to_gpr;
    wire [31:0] preg32_recover_table_to_gpr;
    wire [31:0] preg33_recover_table_to_gpr;
    wire [31:0] preg34_recover_table_to_gpr;
    wire [31:0] preg35_recover_table_to_gpr;
    wire [31:0] preg36_recover_table_to_gpr;
    wire [31:0] preg37_recover_table_to_gpr;
    wire [31:0] preg38_recover_table_to_gpr;
    wire [31:0] preg39_recover_table_to_gpr;
    wire [31:0] preg40_recover_table_to_gpr;
    wire [31:0] preg41_recover_table_to_gpr;
    wire [31:0] preg42_recover_table_to_gpr;
    wire [31:0] preg43_recover_table_to_gpr;
    wire [31:0] preg44_recover_table_to_gpr;
    wire [31:0] preg45_recover_table_to_gpr;
    wire [31:0] preg46_recover_table_to_gpr;
    wire [31:0] preg47_recover_table_to_gpr;
    wire [31:0] preg48_recover_table_to_gpr;
    wire [31:0] preg49_recover_table_to_gpr;
    wire [31:0] preg50_recover_table_to_gpr;
    wire [31:0] preg51_recover_table_to_gpr;
    wire [31:0] preg52_recover_table_to_gpr;
    wire [31:0] preg53_recover_table_to_gpr;
    wire [31:0] preg54_recover_table_to_gpr;
    wire [31:0] preg55_recover_table_to_gpr;
    wire [31:0] preg56_recover_table_to_gpr;
    wire [31:0] preg57_recover_table_to_gpr;
    wire [31:0] preg58_recover_table_to_gpr;
    wire [31:0] preg59_recover_table_to_gpr;
    wire [31:0] preg60_recover_table_to_gpr;
    wire [31:0] preg61_recover_table_to_gpr;
    wire [31:0] preg62_recover_table_to_gpr;
    wire [31:0] preg63_recover_table_to_gpr;
    wire [63:0] gpr0_recover_table;
    wire [63:0] gpr1_recover_table;
    wire [63:0] gpr2_recover_table;
    wire [63:0] gpr3_recover_table;
    wire [63:0] gpr4_recover_table;
    wire [63:0] gpr5_recover_table;
    wire [63:0] gpr6_recover_table;
    wire [63:0] gpr7_recover_table;
    wire [63:0] gpr8_recover_table;
    wire [63:0] gpr9_recover_table;
    wire [63:0] gpr10_recover_table;
    wire [63:0] gpr11_recover_table;
    wire [63:0] gpr12_recover_table;
    wire [63:0] gpr13_recover_table;
    wire [63:0] gpr14_recover_table;
    wire [63:0] gpr15_recover_table;
    wire [63:0] gpr16_recover_table;
    wire [63:0] gpr17_recover_table;
    wire [63:0] gpr18_recover_table;
    wire [63:0] gpr19_recover_table;
    wire [63:0] gpr20_recover_table;
    wire [63:0] gpr21_recover_table;
    wire [63:0] gpr22_recover_table;
    wire [63:0] gpr23_recover_table;
    wire [63:0] gpr24_recover_table;
    wire [63:0] gpr25_recover_table;
    wire [63:0] gpr26_recover_table;
    wire [63:0] gpr27_recover_table;
    wire [63:0] gpr28_recover_table;
    wire [63:0] gpr29_recover_table;
    wire [63:0] gpr30_recover_table;
    wire [63:0] gpr31_recover_table;
    wire [5 :0] gpr0_recover_mapped;
    wire [5 :0] gpr1_recover_mapped;
    wire [5 :0] gpr2_recover_mapped;
    wire [5 :0] gpr3_recover_mapped;
    wire [5 :0] gpr4_recover_mapped;
    wire [5 :0] gpr5_recover_mapped;
    wire [5 :0] gpr6_recover_mapped;
    wire [5 :0] gpr7_recover_mapped;
    wire [5 :0] gpr8_recover_mapped;
    wire [5 :0] gpr9_recover_mapped;
    wire [5 :0] gpr10_recover_mapped;
    wire [5 :0] gpr11_recover_mapped;
    wire [5 :0] gpr12_recover_mapped;
    wire [5 :0] gpr13_recover_mapped;
    wire [5 :0] gpr14_recover_mapped;
    wire [5 :0] gpr15_recover_mapped;
    wire [5 :0] gpr16_recover_mapped;
    wire [5 :0] gpr17_recover_mapped;
    wire [5 :0] gpr18_recover_mapped;
    wire [5 :0] gpr19_recover_mapped;
    wire [5 :0] gpr20_recover_mapped;
    wire [5 :0] gpr21_recover_mapped;
    wire [5 :0] gpr22_recover_mapped;
    wire [5 :0] gpr23_recover_mapped;
    wire [5 :0] gpr24_recover_mapped;
    wire [5 :0] gpr25_recover_mapped;
    wire [5 :0] gpr26_recover_mapped;
    wire [5 :0] gpr27_recover_mapped;
    wire [5 :0] gpr28_recover_mapped;
    wire [5 :0] gpr29_recover_mapped;
    wire [5 :0] gpr30_recover_mapped;
    wire [5 :0] gpr31_recover_mapped;

    // entrys
    assign preg0_release_expand       = 64'b0;
    assign preg0_recover_table_to_gpr = 32'b1;
    assign preg_dealloc[0]            = 1'b0;

    rtu_pst_preg_entry rtu_pst_preg1_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[1]              ),
        .x_alloc_vld                    (preg_alloc_vld[1]                  ),
        .x_release_vld                  (preg_release_vld[1]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[1]              ),
        .x_reset_mapped                 (preg_reset_mapped[1]               ),
        .x_reset_gpr_mapped             (preg1_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg1_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg1_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[1]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg2_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[2]              ),
        .x_alloc_vld                    (preg_alloc_vld[2]                  ),
        .x_release_vld                  (preg_release_vld[2]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[2]              ),
        .x_reset_mapped                 (preg_reset_mapped[2]               ),
        .x_reset_gpr_mapped             (preg2_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg2_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg2_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[2]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg3_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[3]              ),
        .x_alloc_vld                    (preg_alloc_vld[3]                  ),
        .x_release_vld                  (preg_release_vld[3]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[3]              ),
        .x_reset_mapped                 (preg_reset_mapped[3]               ),
        .x_reset_gpr_mapped             (preg3_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg3_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg3_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[3]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg4_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[4]              ),
        .x_alloc_vld                    (preg_alloc_vld[4]                  ),
        .x_release_vld                  (preg_release_vld[4]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[4]              ),
        .x_reset_mapped                 (preg_reset_mapped[4]               ),
        .x_reset_gpr_mapped             (preg4_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg4_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg4_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[4]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg5_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[5]              ),
        .x_alloc_vld                    (preg_alloc_vld[5]                  ),
        .x_release_vld                  (preg_release_vld[5]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[5]              ),
        .x_reset_mapped                 (preg_reset_mapped[5]               ),
        .x_reset_gpr_mapped             (preg5_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg5_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg5_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[5]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg6_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[6]              ),
        .x_alloc_vld                    (preg_alloc_vld[6]                  ),
        .x_release_vld                  (preg_release_vld[6]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[6]              ),
        .x_reset_mapped                 (preg_reset_mapped[6]               ),
        .x_reset_gpr_mapped             (preg6_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg6_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg6_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[6]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg7_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[7]              ),
        .x_alloc_vld                    (preg_alloc_vld[7]                  ),
        .x_release_vld                  (preg_release_vld[7]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[7]              ),
        .x_reset_mapped                 (preg_reset_mapped[7]               ),
        .x_reset_gpr_mapped             (preg7_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg7_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg7_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[7]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg8_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[8]              ),
        .x_alloc_vld                    (preg_alloc_vld[8]                  ),
        .x_release_vld                  (preg_release_vld[8]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[8]              ),
        .x_reset_mapped                 (preg_reset_mapped[8]               ),
        .x_reset_gpr_mapped             (preg8_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg8_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg8_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[8]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg9_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[9]              ),
        .x_alloc_vld                    (preg_alloc_vld[9]                  ),
        .x_release_vld                  (preg_release_vld[9]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[9]              ),
        .x_reset_mapped                 (preg_reset_mapped[9]               ),
        .x_reset_gpr_mapped             (preg9_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg9_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg9_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[9]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg10_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[10]              ),
        .x_alloc_vld                    (preg_alloc_vld[10]                  ),
        .x_release_vld                  (preg_release_vld[10]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[10]              ),
        .x_reset_mapped                 (preg_reset_mapped[10]               ),
        .x_reset_gpr_mapped             (preg10_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg10_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg10_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[10]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg11_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[11]              ),
        .x_alloc_vld                    (preg_alloc_vld[11]                  ),
        .x_release_vld                  (preg_release_vld[11]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[11]              ),
        .x_reset_mapped                 (preg_reset_mapped[11]               ),
        .x_reset_gpr_mapped             (preg11_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg11_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg11_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[11]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg12_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[12]              ),
        .x_alloc_vld                    (preg_alloc_vld[12]                  ),
        .x_release_vld                  (preg_release_vld[12]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[12]              ),
        .x_reset_mapped                 (preg_reset_mapped[12]               ),
        .x_reset_gpr_mapped             (preg12_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg12_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg12_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[12]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg13_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[13]              ),
        .x_alloc_vld                    (preg_alloc_vld[13]                  ),
        .x_release_vld                  (preg_release_vld[13]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[13]              ),
        .x_reset_mapped                 (preg_reset_mapped[13]               ),
        .x_reset_gpr_mapped             (preg13_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg13_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg13_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[13]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg14_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[14]              ),
        .x_alloc_vld                    (preg_alloc_vld[14]                  ),
        .x_release_vld                  (preg_release_vld[14]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[14]              ),
        .x_reset_mapped                 (preg_reset_mapped[14]               ),
        .x_reset_gpr_mapped             (preg14_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg14_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg14_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[14]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg15_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[15]              ),
        .x_alloc_vld                    (preg_alloc_vld[15]                  ),
        .x_release_vld                  (preg_release_vld[15]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[15]              ),
        .x_reset_mapped                 (preg_reset_mapped[15]               ),
        .x_reset_gpr_mapped             (preg15_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg15_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg15_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[15]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg16_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[16]              ),
        .x_alloc_vld                    (preg_alloc_vld[16]                  ),
        .x_release_vld                  (preg_release_vld[16]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[16]              ),
        .x_reset_mapped                 (preg_reset_mapped[16]               ),
        .x_reset_gpr_mapped             (preg16_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg16_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg16_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[16]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg17_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[17]              ),
        .x_alloc_vld                    (preg_alloc_vld[17]                  ),
        .x_release_vld                  (preg_release_vld[17]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[17]              ),
        .x_reset_mapped                 (preg_reset_mapped[17]               ),
        .x_reset_gpr_mapped             (preg17_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg17_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg17_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[17]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg18_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[18]              ),
        .x_alloc_vld                    (preg_alloc_vld[18]                  ),
        .x_release_vld                  (preg_release_vld[18]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[18]              ),
        .x_reset_mapped                 (preg_reset_mapped[18]               ),
        .x_reset_gpr_mapped             (preg18_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg18_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg18_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[18]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg19_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[19]              ),
        .x_alloc_vld                    (preg_alloc_vld[19]                  ),
        .x_release_vld                  (preg_release_vld[19]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[19]              ),
        .x_reset_mapped                 (preg_reset_mapped[19]               ),
        .x_reset_gpr_mapped             (preg19_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg19_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg19_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[19]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg20_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[20]              ),
        .x_alloc_vld                    (preg_alloc_vld[20]                  ),
        .x_release_vld                  (preg_release_vld[20]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[20]              ),
        .x_reset_mapped                 (preg_reset_mapped[20]               ),
        .x_reset_gpr_mapped             (preg20_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg20_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg20_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[20]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg21_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[21]              ),
        .x_alloc_vld                    (preg_alloc_vld[21]                  ),
        .x_release_vld                  (preg_release_vld[21]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[21]              ),
        .x_reset_mapped                 (preg_reset_mapped[21]               ),
        .x_reset_gpr_mapped             (preg21_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg21_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg21_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[21]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg22_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[22]              ),
        .x_alloc_vld                    (preg_alloc_vld[22]                  ),
        .x_release_vld                  (preg_release_vld[22]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[22]              ),
        .x_reset_mapped                 (preg_reset_mapped[22]               ),
        .x_reset_gpr_mapped             (preg22_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg22_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg22_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[22]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg23_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[23]              ),
        .x_alloc_vld                    (preg_alloc_vld[23]                  ),
        .x_release_vld                  (preg_release_vld[23]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[23]              ),
        .x_reset_mapped                 (preg_reset_mapped[23]               ),
        .x_reset_gpr_mapped             (preg23_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg23_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg23_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[23]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg24_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[24]              ),
        .x_alloc_vld                    (preg_alloc_vld[24]                  ),
        .x_release_vld                  (preg_release_vld[24]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[24]              ),
        .x_reset_mapped                 (preg_reset_mapped[24]               ),
        .x_reset_gpr_mapped             (preg24_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg24_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg24_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[24]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg25_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[25]              ),
        .x_alloc_vld                    (preg_alloc_vld[25]                  ),
        .x_release_vld                  (preg_release_vld[25]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[25]              ),
        .x_reset_mapped                 (preg_reset_mapped[25]               ),
        .x_reset_gpr_mapped             (preg25_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg25_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg25_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[25]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg26_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[26]              ),
        .x_alloc_vld                    (preg_alloc_vld[26]                  ),
        .x_release_vld                  (preg_release_vld[26]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[26]              ),
        .x_reset_mapped                 (preg_reset_mapped[26]               ),
        .x_reset_gpr_mapped             (preg26_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg26_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg26_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[26]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg27_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[27]              ),
        .x_alloc_vld                    (preg_alloc_vld[27]                  ),
        .x_release_vld                  (preg_release_vld[27]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[27]              ),
        .x_reset_mapped                 (preg_reset_mapped[27]               ),
        .x_reset_gpr_mapped             (preg27_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg27_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg27_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[27]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg28_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[28]              ),
        .x_alloc_vld                    (preg_alloc_vld[28]                  ),
        .x_release_vld                  (preg_release_vld[28]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[28]              ),
        .x_reset_mapped                 (preg_reset_mapped[28]               ),
        .x_reset_gpr_mapped             (preg28_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg28_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg28_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[28]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg29_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[29]              ),
        .x_alloc_vld                    (preg_alloc_vld[29]                  ),
        .x_release_vld                  (preg_release_vld[29]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[29]              ),
        .x_reset_mapped                 (preg_reset_mapped[29]               ),
        .x_reset_gpr_mapped             (preg29_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg29_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg29_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[29]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg30_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[30]              ),
        .x_alloc_vld                    (preg_alloc_vld[30]                  ),
        .x_release_vld                  (preg_release_vld[30]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[30]              ),
        .x_reset_mapped                 (preg_reset_mapped[30]               ),
        .x_reset_gpr_mapped             (preg30_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg30_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg30_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[30]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg31_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[31]              ),
        .x_alloc_vld                    (preg_alloc_vld[31]                  ),
        .x_release_vld                  (preg_release_vld[31]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[31]              ),
        .x_reset_mapped                 (preg_reset_mapped[31]               ),
        .x_reset_gpr_mapped             (preg31_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg31_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg31_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[31]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg32_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[32]              ),
        .x_alloc_vld                    (preg_alloc_vld[32]                  ),
        .x_release_vld                  (preg_release_vld[32]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[32]              ),
        .x_reset_mapped                 (preg_reset_mapped[32]               ),
        .x_reset_gpr_mapped             (preg32_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg32_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg32_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[32]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg33_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[33]              ),
        .x_alloc_vld                    (preg_alloc_vld[33]                  ),
        .x_release_vld                  (preg_release_vld[33]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[33]              ),
        .x_reset_mapped                 (preg_reset_mapped[33]               ),
        .x_reset_gpr_mapped             (preg33_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg33_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg33_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[33]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg34_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[34]              ),
        .x_alloc_vld                    (preg_alloc_vld[34]                  ),
        .x_release_vld                  (preg_release_vld[34]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[34]              ),
        .x_reset_mapped                 (preg_reset_mapped[34]               ),
        .x_reset_gpr_mapped             (preg34_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg34_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg34_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[34]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg35_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[35]              ),
        .x_alloc_vld                    (preg_alloc_vld[35]                  ),
        .x_release_vld                  (preg_release_vld[35]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[35]              ),
        .x_reset_mapped                 (preg_reset_mapped[35]               ),
        .x_reset_gpr_mapped             (preg35_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg35_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg35_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[35]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg36_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[36]              ),
        .x_alloc_vld                    (preg_alloc_vld[36]                  ),
        .x_release_vld                  (preg_release_vld[36]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[36]              ),
        .x_reset_mapped                 (preg_reset_mapped[36]               ),
        .x_reset_gpr_mapped             (preg36_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg36_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg36_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[36]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg37_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[37]              ),
        .x_alloc_vld                    (preg_alloc_vld[37]                  ),
        .x_release_vld                  (preg_release_vld[37]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[37]              ),
        .x_reset_mapped                 (preg_reset_mapped[37]               ),
        .x_reset_gpr_mapped             (preg37_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg37_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg37_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[37]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg38_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[38]              ),
        .x_alloc_vld                    (preg_alloc_vld[38]                  ),
        .x_release_vld                  (preg_release_vld[38]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[38]              ),
        .x_reset_mapped                 (preg_reset_mapped[38]               ),
        .x_reset_gpr_mapped             (preg38_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg38_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg38_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[38]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg39_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[39]              ),
        .x_alloc_vld                    (preg_alloc_vld[39]                  ),
        .x_release_vld                  (preg_release_vld[39]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[39]              ),
        .x_reset_mapped                 (preg_reset_mapped[39]               ),
        .x_reset_gpr_mapped             (preg39_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg39_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg39_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[39]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg40_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[40]              ),
        .x_alloc_vld                    (preg_alloc_vld[40]                  ),
        .x_release_vld                  (preg_release_vld[40]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[40]              ),
        .x_reset_mapped                 (preg_reset_mapped[40]               ),
        .x_reset_gpr_mapped             (preg40_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg40_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg40_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[40]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg41_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[41]              ),
        .x_alloc_vld                    (preg_alloc_vld[41]                  ),
        .x_release_vld                  (preg_release_vld[41]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[41]              ),
        .x_reset_mapped                 (preg_reset_mapped[41]               ),
        .x_reset_gpr_mapped             (preg41_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg41_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg41_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[41]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg42_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[42]              ),
        .x_alloc_vld                    (preg_alloc_vld[42]                  ),
        .x_release_vld                  (preg_release_vld[42]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[42]              ),
        .x_reset_mapped                 (preg_reset_mapped[42]               ),
        .x_reset_gpr_mapped             (preg42_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg42_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg42_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[42]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg43_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[43]              ),
        .x_alloc_vld                    (preg_alloc_vld[43]                  ),
        .x_release_vld                  (preg_release_vld[43]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[43]              ),
        .x_reset_mapped                 (preg_reset_mapped[43]               ),
        .x_reset_gpr_mapped             (preg43_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg43_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg43_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[43]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg44_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[44]              ),
        .x_alloc_vld                    (preg_alloc_vld[44]                  ),
        .x_release_vld                  (preg_release_vld[44]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[44]              ),
        .x_reset_mapped                 (preg_reset_mapped[44]               ),
        .x_reset_gpr_mapped             (preg44_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg44_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg44_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[44]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg45_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[45]              ),
        .x_alloc_vld                    (preg_alloc_vld[45]                  ),
        .x_release_vld                  (preg_release_vld[45]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[45]              ),
        .x_reset_mapped                 (preg_reset_mapped[45]               ),
        .x_reset_gpr_mapped             (preg45_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg45_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg45_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[45]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg46_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[46]              ),
        .x_alloc_vld                    (preg_alloc_vld[46]                  ),
        .x_release_vld                  (preg_release_vld[46]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[46]              ),
        .x_reset_mapped                 (preg_reset_mapped[46]               ),
        .x_reset_gpr_mapped             (preg46_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg46_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg46_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[46]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg47_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[47]              ),
        .x_alloc_vld                    (preg_alloc_vld[47]                  ),
        .x_release_vld                  (preg_release_vld[47]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[47]              ),
        .x_reset_mapped                 (preg_reset_mapped[47]               ),
        .x_reset_gpr_mapped             (preg47_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg47_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg47_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[47]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg48_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[48]              ),
        .x_alloc_vld                    (preg_alloc_vld[48]                  ),
        .x_release_vld                  (preg_release_vld[48]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[48]              ),
        .x_reset_mapped                 (preg_reset_mapped[48]               ),
        .x_reset_gpr_mapped             (preg48_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg48_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg48_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[48]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg49_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[49]              ),
        .x_alloc_vld                    (preg_alloc_vld[49]                  ),
        .x_release_vld                  (preg_release_vld[49]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[49]              ),
        .x_reset_mapped                 (preg_reset_mapped[49]               ),
        .x_reset_gpr_mapped             (preg49_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg49_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg49_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[49]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg50_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[50]              ),
        .x_alloc_vld                    (preg_alloc_vld[50]                  ),
        .x_release_vld                  (preg_release_vld[50]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[50]              ),
        .x_reset_mapped                 (preg_reset_mapped[50]               ),
        .x_reset_gpr_mapped             (preg50_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg50_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg50_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[50]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg51_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[51]              ),
        .x_alloc_vld                    (preg_alloc_vld[51]                  ),
        .x_release_vld                  (preg_release_vld[51]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[51]              ),
        .x_reset_mapped                 (preg_reset_mapped[51]               ),
        .x_reset_gpr_mapped             (preg51_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg51_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg51_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[51]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg52_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[52]              ),
        .x_alloc_vld                    (preg_alloc_vld[52]                  ),
        .x_release_vld                  (preg_release_vld[52]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[52]              ),
        .x_reset_mapped                 (preg_reset_mapped[52]               ),
        .x_reset_gpr_mapped             (preg52_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg52_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg52_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[52]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg53_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[53]              ),
        .x_alloc_vld                    (preg_alloc_vld[53]                  ),
        .x_release_vld                  (preg_release_vld[53]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[53]              ),
        .x_reset_mapped                 (preg_reset_mapped[53]               ),
        .x_reset_gpr_mapped             (preg53_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg53_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg53_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[53]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg54_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[54]              ),
        .x_alloc_vld                    (preg_alloc_vld[54]                  ),
        .x_release_vld                  (preg_release_vld[54]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[54]              ),
        .x_reset_mapped                 (preg_reset_mapped[54]               ),
        .x_reset_gpr_mapped             (preg54_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg54_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg54_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[54]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg55_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[55]              ),
        .x_alloc_vld                    (preg_alloc_vld[55]                  ),
        .x_release_vld                  (preg_release_vld[55]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[55]              ),
        .x_reset_mapped                 (preg_reset_mapped[55]               ),
        .x_reset_gpr_mapped             (preg55_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg55_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg55_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[55]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg56_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[56]              ),
        .x_alloc_vld                    (preg_alloc_vld[56]                  ),
        .x_release_vld                  (preg_release_vld[56]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[56]              ),
        .x_reset_mapped                 (preg_reset_mapped[56]               ),
        .x_reset_gpr_mapped             (preg56_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg56_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg56_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[56]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg57_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[57]              ),
        .x_alloc_vld                    (preg_alloc_vld[57]                  ),
        .x_release_vld                  (preg_release_vld[57]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[57]              ),
        .x_reset_mapped                 (preg_reset_mapped[57]               ),
        .x_reset_gpr_mapped             (preg57_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg57_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg57_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[57]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg58_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[58]              ),
        .x_alloc_vld                    (preg_alloc_vld[58]                  ),
        .x_release_vld                  (preg_release_vld[58]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[58]              ),
        .x_reset_mapped                 (preg_reset_mapped[58]               ),
        .x_reset_gpr_mapped             (preg58_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg58_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg58_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[58]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg59_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[59]              ),
        .x_alloc_vld                    (preg_alloc_vld[59]                  ),
        .x_release_vld                  (preg_release_vld[59]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[59]              ),
        .x_reset_mapped                 (preg_reset_mapped[59]               ),
        .x_reset_gpr_mapped             (preg59_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg59_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg59_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[59]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg60_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[60]              ),
        .x_alloc_vld                    (preg_alloc_vld[60]                  ),
        .x_release_vld                  (preg_release_vld[60]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[60]              ),
        .x_reset_mapped                 (preg_reset_mapped[60]               ),
        .x_reset_gpr_mapped             (preg60_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg60_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg60_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[60]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg61_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[61]              ),
        .x_alloc_vld                    (preg_alloc_vld[61]                  ),
        .x_release_vld                  (preg_release_vld[61]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[61]              ),
        .x_reset_mapped                 (preg_reset_mapped[61]               ),
        .x_reset_gpr_mapped             (preg61_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg61_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg61_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[61]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg62_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[62]              ),
        .x_alloc_vld                    (preg_alloc_vld[62]                  ),
        .x_release_vld                  (preg_release_vld[62]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[62]              ),
        .x_reset_mapped                 (preg_reset_mapped[62]               ),
        .x_reset_gpr_mapped             (preg62_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg62_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg62_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[62]                    )
    );

    rtu_pst_preg_entry rtu_pst_preg63_entry(
        .clk                            (clk                                    ),
        .rst_clk                        (rst_clk                                ),
        .create_iid                     (idu_rtu_pst_create_iid                 ),
        .create_gpr_index               (idu_rtu_pst_create_gpr_index           ),
        .create_gpr_pre_preg_index      (idu_rtu_pst_create_gpr_pre_preg_index  ),
        .rtu_global_flush               (rtu_global_flush                       ),
        .x_pre_alloc_vld                (preg_pre_alloc_vld[63]              ),
        .x_alloc_vld                    (preg_alloc_vld[63]                  ),
        .x_release_vld                  (preg_release_vld[63]                ),
        .x_inst_retire_iid              (x_inst_retire_iid                      ),
        .x_retire_vld                   (x_retire_vld                           ),
        .x_wb_vld                       (idu_rtu_pst_wb_vld[63]              ),
        .x_reset_mapped                 (preg_reset_mapped[63]               ),
        .x_reset_gpr_mapped             (preg63_reset_gpr_mapped             ),
        .x_pre_preg_release_expand      (preg63_release_expand               ),
        .x_recover_table_preg_to_gpr    (preg63_recover_table_to_gpr         ),
        .x_preg_cur_stats_dealloc       (preg_dealloc[63]                    )
    );

    // pre alloc priority

    assign preg_pre_alloc_priority[0]  = preg_dealloc[0];
    assign preg_pre_alloc_priority[1]  = preg_dealloc[1]  && !preg_dealloc[0];
    assign preg_pre_alloc_priority[2]  = preg_dealloc[2]  && !(|preg_dealloc[1:0]);
    assign preg_pre_alloc_priority[3]  = preg_dealloc[3]  && !(|preg_dealloc[2:0]);
    assign preg_pre_alloc_priority[4]  = preg_dealloc[4]  && !(|preg_dealloc[3:0]);
    assign preg_pre_alloc_priority[5]  = preg_dealloc[5]  && !(|preg_dealloc[4:0]);
    assign preg_pre_alloc_priority[6]  = preg_dealloc[6]  && !(|preg_dealloc[5:0]);
    assign preg_pre_alloc_priority[7]  = preg_dealloc[7]  && !(|preg_dealloc[6:0]);
    assign preg_pre_alloc_priority[8]  = preg_dealloc[8]  && !(|preg_dealloc[7:0]);
    assign preg_pre_alloc_priority[9]  = preg_dealloc[9]  && !(|preg_dealloc[8:0]);
    assign preg_pre_alloc_priority[10] = preg_dealloc[10] && !(|preg_dealloc[9:0]);
    assign preg_pre_alloc_priority[11] = preg_dealloc[11] && !(|preg_dealloc[10:0]);
    assign preg_pre_alloc_priority[12] = preg_dealloc[12] && !(|preg_dealloc[11:0]);
    assign preg_pre_alloc_priority[13] = preg_dealloc[13] && !(|preg_dealloc[12:0]);
    assign preg_pre_alloc_priority[14] = preg_dealloc[14] && !(|preg_dealloc[13:0]);
    assign preg_pre_alloc_priority[15] = preg_dealloc[15] && !(|preg_dealloc[14:0]);
    assign preg_pre_alloc_priority[16] = preg_dealloc[16] && !(|preg_dealloc[15:0]);
    assign preg_pre_alloc_priority[17] = preg_dealloc[17] && !(|preg_dealloc[16:0]);
    assign preg_pre_alloc_priority[18] = preg_dealloc[18] && !(|preg_dealloc[17:0]);
    assign preg_pre_alloc_priority[19] = preg_dealloc[19] && !(|preg_dealloc[18:0]);
    assign preg_pre_alloc_priority[20] = preg_dealloc[20] && !(|preg_dealloc[19:0]);
    assign preg_pre_alloc_priority[21] = preg_dealloc[21] && !(|preg_dealloc[20:0]);
    assign preg_pre_alloc_priority[22] = preg_dealloc[22] && !(|preg_dealloc[21:0]);
    assign preg_pre_alloc_priority[23] = preg_dealloc[23] && !(|preg_dealloc[22:0]);
    assign preg_pre_alloc_priority[24] = preg_dealloc[24] && !(|preg_dealloc[23:0]);
    assign preg_pre_alloc_priority[25] = preg_dealloc[25] && !(|preg_dealloc[24:0]);
    assign preg_pre_alloc_priority[26] = preg_dealloc[26] && !(|preg_dealloc[25:0]);
    assign preg_pre_alloc_priority[27] = preg_dealloc[27] && !(|preg_dealloc[26:0]);
    assign preg_pre_alloc_priority[28] = preg_dealloc[28] && !(|preg_dealloc[27:0]);
    assign preg_pre_alloc_priority[29] = preg_dealloc[29] && !(|preg_dealloc[28:0]);
    assign preg_pre_alloc_priority[30] = preg_dealloc[30] && !(|preg_dealloc[29:0]);
    assign preg_pre_alloc_priority[31] = preg_dealloc[31] && !(|preg_dealloc[30:0]);
    assign preg_pre_alloc_priority[32] = preg_dealloc[32] && !(|preg_dealloc[31:0]);
    assign preg_pre_alloc_priority[33] = preg_dealloc[33] && !(|preg_dealloc[32:0]);
    assign preg_pre_alloc_priority[34] = preg_dealloc[34] && !(|preg_dealloc[33:0]);
    assign preg_pre_alloc_priority[35] = preg_dealloc[35] && !(|preg_dealloc[34:0]);
    assign preg_pre_alloc_priority[36] = preg_dealloc[36] && !(|preg_dealloc[35:0]);
    assign preg_pre_alloc_priority[37] = preg_dealloc[37] && !(|preg_dealloc[36:0]);
    assign preg_pre_alloc_priority[38] = preg_dealloc[38] && !(|preg_dealloc[37:0]);
    assign preg_pre_alloc_priority[39] = preg_dealloc[39] && !(|preg_dealloc[38:0]);
    assign preg_pre_alloc_priority[40] = preg_dealloc[40] && !(|preg_dealloc[39:0]);
    assign preg_pre_alloc_priority[41] = preg_dealloc[41] && !(|preg_dealloc[40:0]);
    assign preg_pre_alloc_priority[42] = preg_dealloc[42] && !(|preg_dealloc[41:0]);
    assign preg_pre_alloc_priority[43] = preg_dealloc[43] && !(|preg_dealloc[42:0]);
    assign preg_pre_alloc_priority[44] = preg_dealloc[44] && !(|preg_dealloc[43:0]);
    assign preg_pre_alloc_priority[45] = preg_dealloc[45] && !(|preg_dealloc[44:0]);
    assign preg_pre_alloc_priority[46] = preg_dealloc[46] && !(|preg_dealloc[45:0]);
    assign preg_pre_alloc_priority[47] = preg_dealloc[47] && !(|preg_dealloc[46:0]);
    assign preg_pre_alloc_priority[48] = preg_dealloc[48] && !(|preg_dealloc[47:0]);
    assign preg_pre_alloc_priority[49] = preg_dealloc[49] && !(|preg_dealloc[48:0]);
    assign preg_pre_alloc_priority[50] = preg_dealloc[50] && !(|preg_dealloc[49:0]);
    assign preg_pre_alloc_priority[51] = preg_dealloc[51] && !(|preg_dealloc[50:0]);
    assign preg_pre_alloc_priority[52] = preg_dealloc[52] && !(|preg_dealloc[51:0]);
    assign preg_pre_alloc_priority[53] = preg_dealloc[53] && !(|preg_dealloc[52:0]);
    assign preg_pre_alloc_priority[54] = preg_dealloc[54] && !(|preg_dealloc[53:0]);
    assign preg_pre_alloc_priority[55] = preg_dealloc[55] && !(|preg_dealloc[54:0]);
    assign preg_pre_alloc_priority[56] = preg_dealloc[56] && !(|preg_dealloc[55:0]);
    assign preg_pre_alloc_priority[57] = preg_dealloc[57] && !(|preg_dealloc[56:0]);
    assign preg_pre_alloc_priority[58] = preg_dealloc[58] && !(|preg_dealloc[57:0]);
    assign preg_pre_alloc_priority[59] = preg_dealloc[59] && !(|preg_dealloc[58:0]);
    assign preg_pre_alloc_priority[60] = preg_dealloc[60] && !(|preg_dealloc[59:0]);
    assign preg_pre_alloc_priority[61] = preg_dealloc[61] && !(|preg_dealloc[60:0]);
    assign preg_pre_alloc_priority[62] = preg_dealloc[62] && !(|preg_dealloc[61:0]);
    assign preg_pre_alloc_priority[63] = preg_dealloc[63] && !(|preg_dealloc[62:0]);

    assign preg_pre_alloc_vld = preg_pre_alloc_priority & {64{alloc_preg_invalid}};

    assign pre_alloc_preg = {6{preg_pre_alloc_priority[0]}}  & 6'd0
                          | {6{preg_pre_alloc_priority[1]}}  & 6'd1
                          | {6{preg_pre_alloc_priority[2]}}  & 6'd2
                          | {6{preg_pre_alloc_priority[3]}}  & 6'd3
                          | {6{preg_pre_alloc_priority[4]}}  & 6'd4
                          | {6{preg_pre_alloc_priority[5]}}  & 6'd5
                          | {6{preg_pre_alloc_priority[6]}}  & 6'd6
                          | {6{preg_pre_alloc_priority[7]}}  & 6'd7
                          | {6{preg_pre_alloc_priority[8]}}  & 6'd8
                          | {6{preg_pre_alloc_priority[9]}}  & 6'd9
                          | {6{preg_pre_alloc_priority[10]}} & 6'd10
                          | {6{preg_pre_alloc_priority[12]}} & 6'd12
                          | {6{preg_pre_alloc_priority[13]}} & 6'd13
                          | {6{preg_pre_alloc_priority[14]}} & 6'd14
                          | {6{preg_pre_alloc_priority[15]}} & 6'd15
                          | {6{preg_pre_alloc_priority[16]}} & 6'd16
                          | {6{preg_pre_alloc_priority[17]}} & 6'd17
                          | {6{preg_pre_alloc_priority[18]}} & 6'd18
                          | {6{preg_pre_alloc_priority[19]}} & 6'd19
                          | {6{preg_pre_alloc_priority[20]}} & 6'd20
                          | {6{preg_pre_alloc_priority[21]}} & 6'd21
                          | {6{preg_pre_alloc_priority[22]}} & 6'd22
                          | {6{preg_pre_alloc_priority[23]}} & 6'd23
                          | {6{preg_pre_alloc_priority[24]}} & 6'd24
                          | {6{preg_pre_alloc_priority[25]}} & 6'd25
                          | {6{preg_pre_alloc_priority[26]}} & 6'd26
                          | {6{preg_pre_alloc_priority[27]}} & 6'd27
                          | {6{preg_pre_alloc_priority[28]}} & 6'd28
                          | {6{preg_pre_alloc_priority[29]}} & 6'd29
                          | {6{preg_pre_alloc_priority[30]}} & 6'd30
                          | {6{preg_pre_alloc_priority[31]}} & 6'd31
                          | {6{preg_pre_alloc_priority[32]}} & 6'd32
                          | {6{preg_pre_alloc_priority[33]}} & 6'd33
                          | {6{preg_pre_alloc_priority[34]}} & 6'd34
                          | {6{preg_pre_alloc_priority[35]}} & 6'd35
                          | {6{preg_pre_alloc_priority[36]}} & 6'd36
                          | {6{preg_pre_alloc_priority[37]}} & 6'd37
                          | {6{preg_pre_alloc_priority[38]}} & 6'd38
                          | {6{preg_pre_alloc_priority[39]}} & 6'd39
                          | {6{preg_pre_alloc_priority[40]}} & 6'd40
                          | {6{preg_pre_alloc_priority[41]}} & 6'd41
                          | {6{preg_pre_alloc_priority[42]}} & 6'd42
                          | {6{preg_pre_alloc_priority[43]}} & 6'd43
                          | {6{preg_pre_alloc_priority[44]}} & 6'd44
                          | {6{preg_pre_alloc_priority[45]}} & 6'd45
                          | {6{preg_pre_alloc_priority[46]}} & 6'd46
                          | {6{preg_pre_alloc_priority[47]}} & 6'd47
                          | {6{preg_pre_alloc_priority[48]}} & 6'd48
                          | {6{preg_pre_alloc_priority[49]}} & 6'd49
                          | {6{preg_pre_alloc_priority[50]}} & 6'd50
                          | {6{preg_pre_alloc_priority[51]}} & 6'd51
                          | {6{preg_pre_alloc_priority[52]}} & 6'd52
                          | {6{preg_pre_alloc_priority[53]}} & 6'd53
                          | {6{preg_pre_alloc_priority[54]}} & 6'd54
                          | {6{preg_pre_alloc_priority[55]}} & 6'd55
                          | {6{preg_pre_alloc_priority[56]}} & 6'd56
                          | {6{preg_pre_alloc_priority[57]}} & 6'd57
                          | {6{preg_pre_alloc_priority[58]}} & 6'd58
                          | {6{preg_pre_alloc_priority[59]}} & 6'd59
                          | {6{preg_pre_alloc_priority[60]}} & 6'd60
                          | {6{preg_pre_alloc_priority[61]}} & 6'd61
                          | {6{preg_pre_alloc_priority[62]}} & 6'd62
                          | {6{preg_pre_alloc_priority[63]}} & 6'd63;

    // alloc sign
    for (genvar i = 0; i < 64; i++)
    begin: preg_alloc_vld_sign
        assign preg_alloc_vld[i] = (idu_rtu_pst_create_preg_index == i) && idu_rtu_pst_create_vld;
    end

    // release sign
    for (genvar i = 0; i < 64; i++)
    begin: preg_release_vld_sign
        assign preg_release_vld[i] = preg0_release_expand[i]
                                   | preg1_release_expand[i]
                                   | preg2_release_expand[i]
                                   | preg3_release_expand[i]
                                   | preg4_release_expand[i]
                                   | preg5_release_expand[i]
                                   | preg6_release_expand[i]
                                   | preg7_release_expand[i]
                                   | preg8_release_expand[i]
                                   | preg9_release_expand[i]
                                   | preg10_release_expand[i]
                                   | preg11_release_expand[i]
                                   | preg12_release_expand[i]
                                   | preg13_release_expand[i]
                                   | preg14_release_expand[i]
                                   | preg15_release_expand[i]
                                   | preg16_release_expand[i]
                                   | preg17_release_expand[i]
                                   | preg18_release_expand[i]
                                   | preg19_release_expand[i]
                                   | preg20_release_expand[i]
                                   | preg21_release_expand[i]
                                   | preg22_release_expand[i]
                                   | preg23_release_expand[i]
                                   | preg24_release_expand[i]
                                   | preg25_release_expand[i]
                                   | preg26_release_expand[i]
                                   | preg27_release_expand[i]
                                   | preg28_release_expand[i]
                                   | preg29_release_expand[i]
                                   | preg30_release_expand[i]
                                   | preg31_release_expand[i]
                                   | preg32_release_expand[i]
                                   | preg33_release_expand[i]
                                   | preg34_release_expand[i]
                                   | preg35_release_expand[i]
                                   | preg36_release_expand[i]
                                   | preg37_release_expand[i]
                                   | preg38_release_expand[i]
                                   | preg39_release_expand[i]
                                   | preg40_release_expand[i]
                                   | preg41_release_expand[i]
                                   | preg42_release_expand[i]
                                   | preg43_release_expand[i]
                                   | preg44_release_expand[i]
                                   | preg45_release_expand[i]
                                   | preg46_release_expand[i]
                                   | preg47_release_expand[i]
                                   | preg48_release_expand[i]
                                   | preg49_release_expand[i]
                                   | preg50_release_expand[i]
                                   | preg51_release_expand[i]
                                   | preg52_release_expand[i]
                                   | preg53_release_expand[i]
                                   | preg54_release_expand[i]
                                   | preg55_release_expand[i]
                                   | preg56_release_expand[i]
                                   | preg57_release_expand[i]
                                   | preg58_release_expand[i]
                                   | preg59_release_expand[i]
                                   | preg60_release_expand[i]
                                   | preg61_release_expand[i]
                                   | preg62_release_expand[i]
                                   | preg63_release_expand[i];
    end

    // reset vector
    assign preg_reset_mapped = 64'h00000000_ffffffff;
    // assign preg0_reset_gpr_mapped  = 5'd0;
    assign preg1_reset_gpr_mapped  = 5'd1;
    assign preg2_reset_gpr_mapped  = 5'd2;
    assign preg3_reset_gpr_mapped  = 5'd3;
    assign preg4_reset_gpr_mapped  = 5'd4;
    assign preg5_reset_gpr_mapped  = 5'd5;
    assign preg6_reset_gpr_mapped  = 5'd6;
    assign preg7_reset_gpr_mapped  = 5'd7;
    assign preg8_reset_gpr_mapped  = 5'd8;
    assign preg9_reset_gpr_mapped  = 5'd9;
    assign preg10_reset_gpr_mapped = 5'd10;
    assign preg11_reset_gpr_mapped = 5'd11;
    assign preg12_reset_gpr_mapped = 5'd12;
    assign preg13_reset_gpr_mapped = 5'd13;
    assign preg14_reset_gpr_mapped = 5'd14;
    assign preg15_reset_gpr_mapped = 5'd15;
    assign preg16_reset_gpr_mapped = 5'd16;
    assign preg17_reset_gpr_mapped = 5'd17;
    assign preg18_reset_gpr_mapped = 5'd18;
    assign preg19_reset_gpr_mapped = 5'd19;
    assign preg20_reset_gpr_mapped = 5'd20;
    assign preg21_reset_gpr_mapped = 5'd21;
    assign preg22_reset_gpr_mapped = 5'd22;
    assign preg23_reset_gpr_mapped = 5'd23;
    assign preg24_reset_gpr_mapped = 5'd24;
    assign preg25_reset_gpr_mapped = 5'd25;
    assign preg26_reset_gpr_mapped = 5'd26;
    assign preg27_reset_gpr_mapped = 5'd27;
    assign preg28_reset_gpr_mapped = 5'd28;
    assign preg29_reset_gpr_mapped = 5'd29;
    assign preg30_reset_gpr_mapped = 5'd30;
    assign preg31_reset_gpr_mapped = 5'd31;
    assign preg32_reset_gpr_mapped = 5'd0;
    assign preg33_reset_gpr_mapped = 5'd0;
    assign preg34_reset_gpr_mapped = 5'd0;
    assign preg35_reset_gpr_mapped = 5'd0;
    assign preg36_reset_gpr_mapped = 5'd0;
    assign preg37_reset_gpr_mapped = 5'd0;
    assign preg38_reset_gpr_mapped = 5'd0;
    assign preg39_reset_gpr_mapped = 5'd0;
    assign preg40_reset_gpr_mapped = 5'd0;
    assign preg41_reset_gpr_mapped = 5'd0;
    assign preg42_reset_gpr_mapped = 5'd0;
    assign preg43_reset_gpr_mapped = 5'd0;
    assign preg44_reset_gpr_mapped = 5'd0;
    assign preg45_reset_gpr_mapped = 5'd0;
    assign preg46_reset_gpr_mapped = 5'd0;
    assign preg47_reset_gpr_mapped = 5'd0;
    assign preg48_reset_gpr_mapped = 5'd0;
    assign preg49_reset_gpr_mapped = 5'd0;
    assign preg50_reset_gpr_mapped = 5'd0;
    assign preg51_reset_gpr_mapped = 5'd0;
    assign preg52_reset_gpr_mapped = 5'd0;
    assign preg53_reset_gpr_mapped = 5'd0;
    assign preg54_reset_gpr_mapped = 5'd0;
    assign preg55_reset_gpr_mapped = 5'd0;
    assign preg56_reset_gpr_mapped = 5'd0;
    assign preg57_reset_gpr_mapped = 5'd0;
    assign preg58_reset_gpr_mapped = 5'd0;
    assign preg59_reset_gpr_mapped = 5'd0;
    assign preg60_reset_gpr_mapped = 5'd0;
    assign preg61_reset_gpr_mapped = 5'd0;
    assign preg62_reset_gpr_mapped = 5'd0;
    assign preg63_reset_gpr_mapped = 5'd0;

    // recover table
    assign gpr0_recover_table = {preg63_recover_table_to_gpr[0], preg62_recover_table_to_gpr[0], preg61_recover_table_to_gpr[0], preg60_recover_table_to_gpr[0],
                                 preg59_recover_table_to_gpr[0], preg58_recover_table_to_gpr[0], preg57_recover_table_to_gpr[0], preg56_recover_table_to_gpr[0],
                                 preg55_recover_table_to_gpr[0], preg54_recover_table_to_gpr[0], preg53_recover_table_to_gpr[0], preg52_recover_table_to_gpr[0],
                                 preg51_recover_table_to_gpr[0], preg50_recover_table_to_gpr[0], preg49_recover_table_to_gpr[0], preg48_recover_table_to_gpr[0],
                                 preg47_recover_table_to_gpr[0], preg46_recover_table_to_gpr[0], preg45_recover_table_to_gpr[0], preg44_recover_table_to_gpr[0],
                                 preg43_recover_table_to_gpr[0], preg42_recover_table_to_gpr[0], preg41_recover_table_to_gpr[0], preg40_recover_table_to_gpr[0],
                                 preg39_recover_table_to_gpr[0], preg38_recover_table_to_gpr[0], preg37_recover_table_to_gpr[0], preg36_recover_table_to_gpr[0],
                                 preg35_recover_table_to_gpr[0], preg34_recover_table_to_gpr[0], preg33_recover_table_to_gpr[0], preg32_recover_table_to_gpr[0],
                                 preg31_recover_table_to_gpr[0], preg30_recover_table_to_gpr[0], preg29_recover_table_to_gpr[0], preg28_recover_table_to_gpr[0],
                                 preg27_recover_table_to_gpr[0], preg26_recover_table_to_gpr[0], preg25_recover_table_to_gpr[0], preg24_recover_table_to_gpr[0],
                                 preg23_recover_table_to_gpr[0], preg22_recover_table_to_gpr[0], preg21_recover_table_to_gpr[0], preg20_recover_table_to_gpr[0],
                                 preg19_recover_table_to_gpr[0], preg18_recover_table_to_gpr[0], preg17_recover_table_to_gpr[0], preg16_recover_table_to_gpr[0],
                                 preg15_recover_table_to_gpr[0], preg14_recover_table_to_gpr[0], preg13_recover_table_to_gpr[0], preg12_recover_table_to_gpr[0],
                                 preg11_recover_table_to_gpr[0], preg10_recover_table_to_gpr[0], preg9_recover_table_to_gpr[0],  preg8_recover_table_to_gpr[0] ,
                                 preg7_recover_table_to_gpr[0],  preg6_recover_table_to_gpr[0],  preg5_recover_table_to_gpr[0],  preg4_recover_table_to_gpr[0] ,
                                 preg3_recover_table_to_gpr[0],  preg2_recover_table_to_gpr[0],  preg1_recover_table_to_gpr[0],  preg0_recover_table_to_gpr[0]};
    assign gpr1_recover_table = {preg63_recover_table_to_gpr[1], preg62_recover_table_to_gpr[1], preg61_recover_table_to_gpr[1], preg60_recover_table_to_gpr[1],
                                 preg59_recover_table_to_gpr[1], preg58_recover_table_to_gpr[1], preg57_recover_table_to_gpr[1], preg56_recover_table_to_gpr[1],
                                 preg55_recover_table_to_gpr[1], preg54_recover_table_to_gpr[1], preg53_recover_table_to_gpr[1], preg52_recover_table_to_gpr[1],
                                 preg51_recover_table_to_gpr[1], preg50_recover_table_to_gpr[1], preg49_recover_table_to_gpr[1], preg48_recover_table_to_gpr[1],
                                 preg47_recover_table_to_gpr[1], preg46_recover_table_to_gpr[1], preg45_recover_table_to_gpr[1], preg44_recover_table_to_gpr[1],
                                 preg43_recover_table_to_gpr[1], preg42_recover_table_to_gpr[1], preg41_recover_table_to_gpr[1], preg40_recover_table_to_gpr[1],
                                 preg39_recover_table_to_gpr[1], preg38_recover_table_to_gpr[1], preg37_recover_table_to_gpr[1], preg36_recover_table_to_gpr[1],
                                 preg35_recover_table_to_gpr[1], preg34_recover_table_to_gpr[1], preg33_recover_table_to_gpr[1], preg32_recover_table_to_gpr[1],
                                 preg31_recover_table_to_gpr[1], preg30_recover_table_to_gpr[1], preg29_recover_table_to_gpr[1], preg28_recover_table_to_gpr[1],
                                 preg27_recover_table_to_gpr[1], preg26_recover_table_to_gpr[1], preg25_recover_table_to_gpr[1], preg24_recover_table_to_gpr[1],
                                 preg23_recover_table_to_gpr[1], preg22_recover_table_to_gpr[1], preg21_recover_table_to_gpr[1], preg20_recover_table_to_gpr[1],
                                 preg19_recover_table_to_gpr[1], preg18_recover_table_to_gpr[1], preg17_recover_table_to_gpr[1], preg16_recover_table_to_gpr[1],
                                 preg15_recover_table_to_gpr[1], preg14_recover_table_to_gpr[1], preg13_recover_table_to_gpr[1], preg12_recover_table_to_gpr[1],
                                 preg11_recover_table_to_gpr[1], preg10_recover_table_to_gpr[1], preg9_recover_table_to_gpr[1],  preg8_recover_table_to_gpr[1] ,
                                 preg7_recover_table_to_gpr[1],  preg6_recover_table_to_gpr[1],  preg5_recover_table_to_gpr[1],  preg4_recover_table_to_gpr[1] ,
                                 preg3_recover_table_to_gpr[1],  preg2_recover_table_to_gpr[1],  preg1_recover_table_to_gpr[1],  preg0_recover_table_to_gpr[1]};
    assign gpr2_recover_table = {preg63_recover_table_to_gpr[2], preg62_recover_table_to_gpr[2], preg61_recover_table_to_gpr[2], preg60_recover_table_to_gpr[2],
                                 preg59_recover_table_to_gpr[2], preg58_recover_table_to_gpr[2], preg57_recover_table_to_gpr[2], preg56_recover_table_to_gpr[2],
                                 preg55_recover_table_to_gpr[2], preg54_recover_table_to_gpr[2], preg53_recover_table_to_gpr[2], preg52_recover_table_to_gpr[2],
                                 preg51_recover_table_to_gpr[2], preg50_recover_table_to_gpr[2], preg49_recover_table_to_gpr[2], preg48_recover_table_to_gpr[2],
                                 preg47_recover_table_to_gpr[2], preg46_recover_table_to_gpr[2], preg45_recover_table_to_gpr[2], preg44_recover_table_to_gpr[2],
                                 preg43_recover_table_to_gpr[2], preg42_recover_table_to_gpr[2], preg41_recover_table_to_gpr[2], preg40_recover_table_to_gpr[2],
                                 preg39_recover_table_to_gpr[2], preg38_recover_table_to_gpr[2], preg37_recover_table_to_gpr[2], preg36_recover_table_to_gpr[2],
                                 preg35_recover_table_to_gpr[2], preg34_recover_table_to_gpr[2], preg33_recover_table_to_gpr[2], preg32_recover_table_to_gpr[2],
                                 preg31_recover_table_to_gpr[2], preg30_recover_table_to_gpr[2], preg29_recover_table_to_gpr[2], preg28_recover_table_to_gpr[2],
                                 preg27_recover_table_to_gpr[2], preg26_recover_table_to_gpr[2], preg25_recover_table_to_gpr[2], preg24_recover_table_to_gpr[2],
                                 preg23_recover_table_to_gpr[2], preg22_recover_table_to_gpr[2], preg21_recover_table_to_gpr[2], preg20_recover_table_to_gpr[2],
                                 preg19_recover_table_to_gpr[2], preg18_recover_table_to_gpr[2], preg17_recover_table_to_gpr[2], preg16_recover_table_to_gpr[2],
                                 preg15_recover_table_to_gpr[2], preg14_recover_table_to_gpr[2], preg13_recover_table_to_gpr[2], preg12_recover_table_to_gpr[2],
                                 preg11_recover_table_to_gpr[2], preg10_recover_table_to_gpr[2], preg9_recover_table_to_gpr[2],  preg8_recover_table_to_gpr[2] ,
                                 preg7_recover_table_to_gpr[2],  preg6_recover_table_to_gpr[2],  preg5_recover_table_to_gpr[2],  preg4_recover_table_to_gpr[2] ,
                                 preg3_recover_table_to_gpr[2],  preg2_recover_table_to_gpr[2],  preg1_recover_table_to_gpr[2],  preg0_recover_table_to_gpr[2]};
    assign gpr3_recover_table = {preg63_recover_table_to_gpr[3], preg62_recover_table_to_gpr[3], preg61_recover_table_to_gpr[3], preg60_recover_table_to_gpr[3],
                                 preg59_recover_table_to_gpr[3], preg58_recover_table_to_gpr[3], preg57_recover_table_to_gpr[3], preg56_recover_table_to_gpr[3],
                                 preg55_recover_table_to_gpr[3], preg54_recover_table_to_gpr[3], preg53_recover_table_to_gpr[3], preg52_recover_table_to_gpr[3],
                                 preg51_recover_table_to_gpr[3], preg50_recover_table_to_gpr[3], preg49_recover_table_to_gpr[3], preg48_recover_table_to_gpr[3],
                                 preg47_recover_table_to_gpr[3], preg46_recover_table_to_gpr[3], preg45_recover_table_to_gpr[3], preg44_recover_table_to_gpr[3],
                                 preg43_recover_table_to_gpr[3], preg42_recover_table_to_gpr[3], preg41_recover_table_to_gpr[3], preg40_recover_table_to_gpr[3],
                                 preg39_recover_table_to_gpr[3], preg38_recover_table_to_gpr[3], preg37_recover_table_to_gpr[3], preg36_recover_table_to_gpr[3],
                                 preg35_recover_table_to_gpr[3], preg34_recover_table_to_gpr[3], preg33_recover_table_to_gpr[3], preg32_recover_table_to_gpr[3],
                                 preg31_recover_table_to_gpr[3], preg30_recover_table_to_gpr[3], preg29_recover_table_to_gpr[3], preg28_recover_table_to_gpr[3],
                                 preg27_recover_table_to_gpr[3], preg26_recover_table_to_gpr[3], preg25_recover_table_to_gpr[3], preg24_recover_table_to_gpr[3],
                                 preg23_recover_table_to_gpr[3], preg22_recover_table_to_gpr[3], preg21_recover_table_to_gpr[3], preg20_recover_table_to_gpr[3],
                                 preg19_recover_table_to_gpr[3], preg18_recover_table_to_gpr[3], preg17_recover_table_to_gpr[3], preg16_recover_table_to_gpr[3],
                                 preg15_recover_table_to_gpr[3], preg14_recover_table_to_gpr[3], preg13_recover_table_to_gpr[3], preg12_recover_table_to_gpr[3],
                                 preg11_recover_table_to_gpr[3], preg10_recover_table_to_gpr[3], preg9_recover_table_to_gpr[3],  preg8_recover_table_to_gpr[3] ,
                                 preg7_recover_table_to_gpr[3],  preg6_recover_table_to_gpr[3],  preg5_recover_table_to_gpr[3],  preg4_recover_table_to_gpr[3] ,
                                 preg3_recover_table_to_gpr[3],  preg2_recover_table_to_gpr[3],  preg1_recover_table_to_gpr[3],  preg0_recover_table_to_gpr[3]};
    assign gpr4_recover_table = {preg63_recover_table_to_gpr[4], preg62_recover_table_to_gpr[4], preg61_recover_table_to_gpr[4], preg60_recover_table_to_gpr[4],
                                 preg59_recover_table_to_gpr[4], preg58_recover_table_to_gpr[4], preg57_recover_table_to_gpr[4], preg56_recover_table_to_gpr[4],
                                 preg55_recover_table_to_gpr[4], preg54_recover_table_to_gpr[4], preg53_recover_table_to_gpr[4], preg52_recover_table_to_gpr[4],
                                 preg51_recover_table_to_gpr[4], preg50_recover_table_to_gpr[4], preg49_recover_table_to_gpr[4], preg48_recover_table_to_gpr[4],
                                 preg47_recover_table_to_gpr[4], preg46_recover_table_to_gpr[4], preg45_recover_table_to_gpr[4], preg44_recover_table_to_gpr[4],
                                 preg43_recover_table_to_gpr[4], preg42_recover_table_to_gpr[4], preg41_recover_table_to_gpr[4], preg40_recover_table_to_gpr[4],
                                 preg39_recover_table_to_gpr[4], preg38_recover_table_to_gpr[4], preg37_recover_table_to_gpr[4], preg36_recover_table_to_gpr[4],
                                 preg35_recover_table_to_gpr[4], preg34_recover_table_to_gpr[4], preg33_recover_table_to_gpr[4], preg32_recover_table_to_gpr[4],
                                 preg31_recover_table_to_gpr[4], preg30_recover_table_to_gpr[4], preg29_recover_table_to_gpr[4], preg28_recover_table_to_gpr[4],
                                 preg27_recover_table_to_gpr[4], preg26_recover_table_to_gpr[4], preg25_recover_table_to_gpr[4], preg24_recover_table_to_gpr[4],
                                 preg23_recover_table_to_gpr[4], preg22_recover_table_to_gpr[4], preg21_recover_table_to_gpr[4], preg20_recover_table_to_gpr[4],
                                 preg19_recover_table_to_gpr[4], preg18_recover_table_to_gpr[4], preg17_recover_table_to_gpr[4], preg16_recover_table_to_gpr[4],
                                 preg15_recover_table_to_gpr[4], preg14_recover_table_to_gpr[4], preg13_recover_table_to_gpr[4], preg12_recover_table_to_gpr[4],
                                 preg11_recover_table_to_gpr[4], preg10_recover_table_to_gpr[4], preg9_recover_table_to_gpr[4],  preg8_recover_table_to_gpr[4] ,
                                 preg7_recover_table_to_gpr[4],  preg6_recover_table_to_gpr[4],  preg5_recover_table_to_gpr[4],  preg4_recover_table_to_gpr[4] ,
                                 preg3_recover_table_to_gpr[4],  preg2_recover_table_to_gpr[4],  preg1_recover_table_to_gpr[4],  preg0_recover_table_to_gpr[4]};
    assign gpr5_recover_table = {preg63_recover_table_to_gpr[5], preg62_recover_table_to_gpr[5], preg61_recover_table_to_gpr[5], preg60_recover_table_to_gpr[5],
                                 preg59_recover_table_to_gpr[5], preg58_recover_table_to_gpr[5], preg57_recover_table_to_gpr[5], preg56_recover_table_to_gpr[5],
                                 preg55_recover_table_to_gpr[5], preg54_recover_table_to_gpr[5], preg53_recover_table_to_gpr[5], preg52_recover_table_to_gpr[5],
                                 preg51_recover_table_to_gpr[5], preg50_recover_table_to_gpr[5], preg49_recover_table_to_gpr[5], preg48_recover_table_to_gpr[5],
                                 preg47_recover_table_to_gpr[5], preg46_recover_table_to_gpr[5], preg45_recover_table_to_gpr[5], preg44_recover_table_to_gpr[5],
                                 preg43_recover_table_to_gpr[5], preg42_recover_table_to_gpr[5], preg41_recover_table_to_gpr[5], preg40_recover_table_to_gpr[5],
                                 preg39_recover_table_to_gpr[5], preg38_recover_table_to_gpr[5], preg37_recover_table_to_gpr[5], preg36_recover_table_to_gpr[5],
                                 preg35_recover_table_to_gpr[5], preg34_recover_table_to_gpr[5], preg33_recover_table_to_gpr[5], preg32_recover_table_to_gpr[5],
                                 preg31_recover_table_to_gpr[5], preg30_recover_table_to_gpr[5], preg29_recover_table_to_gpr[5], preg28_recover_table_to_gpr[5],
                                 preg27_recover_table_to_gpr[5], preg26_recover_table_to_gpr[5], preg25_recover_table_to_gpr[5], preg24_recover_table_to_gpr[5],
                                 preg23_recover_table_to_gpr[5], preg22_recover_table_to_gpr[5], preg21_recover_table_to_gpr[5], preg20_recover_table_to_gpr[5],
                                 preg19_recover_table_to_gpr[5], preg18_recover_table_to_gpr[5], preg17_recover_table_to_gpr[5], preg16_recover_table_to_gpr[5],
                                 preg15_recover_table_to_gpr[5], preg14_recover_table_to_gpr[5], preg13_recover_table_to_gpr[5], preg12_recover_table_to_gpr[5],
                                 preg11_recover_table_to_gpr[5], preg10_recover_table_to_gpr[5], preg9_recover_table_to_gpr[5],  preg8_recover_table_to_gpr[5] ,
                                 preg7_recover_table_to_gpr[5],  preg6_recover_table_to_gpr[5],  preg5_recover_table_to_gpr[5],  preg4_recover_table_to_gpr[5] ,
                                 preg3_recover_table_to_gpr[5],  preg2_recover_table_to_gpr[5],  preg1_recover_table_to_gpr[5],  preg0_recover_table_to_gpr[5]};
    assign gpr6_recover_table = {preg63_recover_table_to_gpr[6], preg62_recover_table_to_gpr[6], preg61_recover_table_to_gpr[6], preg60_recover_table_to_gpr[6],
                                 preg59_recover_table_to_gpr[6], preg58_recover_table_to_gpr[6], preg57_recover_table_to_gpr[6], preg56_recover_table_to_gpr[6],
                                 preg55_recover_table_to_gpr[6], preg54_recover_table_to_gpr[6], preg53_recover_table_to_gpr[6], preg52_recover_table_to_gpr[6],
                                 preg51_recover_table_to_gpr[6], preg50_recover_table_to_gpr[6], preg49_recover_table_to_gpr[6], preg48_recover_table_to_gpr[6],
                                 preg47_recover_table_to_gpr[6], preg46_recover_table_to_gpr[6], preg45_recover_table_to_gpr[6], preg44_recover_table_to_gpr[6],
                                 preg43_recover_table_to_gpr[6], preg42_recover_table_to_gpr[6], preg41_recover_table_to_gpr[6], preg40_recover_table_to_gpr[6],
                                 preg39_recover_table_to_gpr[6], preg38_recover_table_to_gpr[6], preg37_recover_table_to_gpr[6], preg36_recover_table_to_gpr[6],
                                 preg35_recover_table_to_gpr[6], preg34_recover_table_to_gpr[6], preg33_recover_table_to_gpr[6], preg32_recover_table_to_gpr[6],
                                 preg31_recover_table_to_gpr[6], preg30_recover_table_to_gpr[6], preg29_recover_table_to_gpr[6], preg28_recover_table_to_gpr[6],
                                 preg27_recover_table_to_gpr[6], preg26_recover_table_to_gpr[6], preg25_recover_table_to_gpr[6], preg24_recover_table_to_gpr[6],
                                 preg23_recover_table_to_gpr[6], preg22_recover_table_to_gpr[6], preg21_recover_table_to_gpr[6], preg20_recover_table_to_gpr[6],
                                 preg19_recover_table_to_gpr[6], preg18_recover_table_to_gpr[6], preg17_recover_table_to_gpr[6], preg16_recover_table_to_gpr[6],
                                 preg15_recover_table_to_gpr[6], preg14_recover_table_to_gpr[6], preg13_recover_table_to_gpr[6], preg12_recover_table_to_gpr[6],
                                 preg11_recover_table_to_gpr[6], preg10_recover_table_to_gpr[6], preg9_recover_table_to_gpr[6],  preg8_recover_table_to_gpr[6] ,
                                 preg7_recover_table_to_gpr[6],  preg6_recover_table_to_gpr[6],  preg5_recover_table_to_gpr[6],  preg4_recover_table_to_gpr[6] ,
                                 preg3_recover_table_to_gpr[6],  preg2_recover_table_to_gpr[6],  preg1_recover_table_to_gpr[6],  preg0_recover_table_to_gpr[6]};
    assign gpr7_recover_table = {preg63_recover_table_to_gpr[7], preg62_recover_table_to_gpr[7], preg61_recover_table_to_gpr[7], preg60_recover_table_to_gpr[7],
                                 preg59_recover_table_to_gpr[7], preg58_recover_table_to_gpr[7], preg57_recover_table_to_gpr[7], preg56_recover_table_to_gpr[7],
                                 preg55_recover_table_to_gpr[7], preg54_recover_table_to_gpr[7], preg53_recover_table_to_gpr[7], preg52_recover_table_to_gpr[7],
                                 preg51_recover_table_to_gpr[7], preg50_recover_table_to_gpr[7], preg49_recover_table_to_gpr[7], preg48_recover_table_to_gpr[7],
                                 preg47_recover_table_to_gpr[7], preg46_recover_table_to_gpr[7], preg45_recover_table_to_gpr[7], preg44_recover_table_to_gpr[7],
                                 preg43_recover_table_to_gpr[7], preg42_recover_table_to_gpr[7], preg41_recover_table_to_gpr[7], preg40_recover_table_to_gpr[7],
                                 preg39_recover_table_to_gpr[7], preg38_recover_table_to_gpr[7], preg37_recover_table_to_gpr[7], preg36_recover_table_to_gpr[7],
                                 preg35_recover_table_to_gpr[7], preg34_recover_table_to_gpr[7], preg33_recover_table_to_gpr[7], preg32_recover_table_to_gpr[7],
                                 preg31_recover_table_to_gpr[7], preg30_recover_table_to_gpr[7], preg29_recover_table_to_gpr[7], preg28_recover_table_to_gpr[7],
                                 preg27_recover_table_to_gpr[7], preg26_recover_table_to_gpr[7], preg25_recover_table_to_gpr[7], preg24_recover_table_to_gpr[7],
                                 preg23_recover_table_to_gpr[7], preg22_recover_table_to_gpr[7], preg21_recover_table_to_gpr[7], preg20_recover_table_to_gpr[7],
                                 preg19_recover_table_to_gpr[7], preg18_recover_table_to_gpr[7], preg17_recover_table_to_gpr[7], preg16_recover_table_to_gpr[7],
                                 preg15_recover_table_to_gpr[7], preg14_recover_table_to_gpr[7], preg13_recover_table_to_gpr[7], preg12_recover_table_to_gpr[7],
                                 preg11_recover_table_to_gpr[7], preg10_recover_table_to_gpr[7], preg9_recover_table_to_gpr[7],  preg8_recover_table_to_gpr[7] ,
                                 preg7_recover_table_to_gpr[7],  preg6_recover_table_to_gpr[7],  preg5_recover_table_to_gpr[7],  preg4_recover_table_to_gpr[7] ,
                                 preg3_recover_table_to_gpr[7],  preg2_recover_table_to_gpr[7],  preg1_recover_table_to_gpr[7],  preg0_recover_table_to_gpr[7]};
    assign gpr8_recover_table = {preg63_recover_table_to_gpr[8], preg62_recover_table_to_gpr[8], preg61_recover_table_to_gpr[8], preg60_recover_table_to_gpr[8],
                                 preg59_recover_table_to_gpr[8], preg58_recover_table_to_gpr[8], preg57_recover_table_to_gpr[8], preg56_recover_table_to_gpr[8],
                                 preg55_recover_table_to_gpr[8], preg54_recover_table_to_gpr[8], preg53_recover_table_to_gpr[8], preg52_recover_table_to_gpr[8],
                                 preg51_recover_table_to_gpr[8], preg50_recover_table_to_gpr[8], preg49_recover_table_to_gpr[8], preg48_recover_table_to_gpr[8],
                                 preg47_recover_table_to_gpr[8], preg46_recover_table_to_gpr[8], preg45_recover_table_to_gpr[8], preg44_recover_table_to_gpr[8],
                                 preg43_recover_table_to_gpr[8], preg42_recover_table_to_gpr[8], preg41_recover_table_to_gpr[8], preg40_recover_table_to_gpr[8],
                                 preg39_recover_table_to_gpr[8], preg38_recover_table_to_gpr[8], preg37_recover_table_to_gpr[8], preg36_recover_table_to_gpr[8],
                                 preg35_recover_table_to_gpr[8], preg34_recover_table_to_gpr[8], preg33_recover_table_to_gpr[8], preg32_recover_table_to_gpr[8],
                                 preg31_recover_table_to_gpr[8], preg30_recover_table_to_gpr[8], preg29_recover_table_to_gpr[8], preg28_recover_table_to_gpr[8],
                                 preg27_recover_table_to_gpr[8], preg26_recover_table_to_gpr[8], preg25_recover_table_to_gpr[8], preg24_recover_table_to_gpr[8],
                                 preg23_recover_table_to_gpr[8], preg22_recover_table_to_gpr[8], preg21_recover_table_to_gpr[8], preg20_recover_table_to_gpr[8],
                                 preg19_recover_table_to_gpr[8], preg18_recover_table_to_gpr[8], preg17_recover_table_to_gpr[8], preg16_recover_table_to_gpr[8],
                                 preg15_recover_table_to_gpr[8], preg14_recover_table_to_gpr[8], preg13_recover_table_to_gpr[8], preg12_recover_table_to_gpr[8],
                                 preg11_recover_table_to_gpr[8], preg10_recover_table_to_gpr[8], preg9_recover_table_to_gpr[8],  preg8_recover_table_to_gpr[8] ,
                                 preg7_recover_table_to_gpr[8],  preg6_recover_table_to_gpr[8],  preg5_recover_table_to_gpr[8],  preg4_recover_table_to_gpr[8] ,
                                 preg3_recover_table_to_gpr[8],  preg2_recover_table_to_gpr[8],  preg1_recover_table_to_gpr[8],  preg0_recover_table_to_gpr[8]};
    assign gpr9_recover_table = {preg63_recover_table_to_gpr[9], preg62_recover_table_to_gpr[9], preg61_recover_table_to_gpr[9], preg60_recover_table_to_gpr[9],
                                 preg59_recover_table_to_gpr[9], preg58_recover_table_to_gpr[9], preg57_recover_table_to_gpr[9], preg56_recover_table_to_gpr[9],
                                 preg55_recover_table_to_gpr[9], preg54_recover_table_to_gpr[9], preg53_recover_table_to_gpr[9], preg52_recover_table_to_gpr[9],
                                 preg51_recover_table_to_gpr[9], preg50_recover_table_to_gpr[9], preg49_recover_table_to_gpr[9], preg48_recover_table_to_gpr[9],
                                 preg47_recover_table_to_gpr[9], preg46_recover_table_to_gpr[9], preg45_recover_table_to_gpr[9], preg44_recover_table_to_gpr[9],
                                 preg43_recover_table_to_gpr[9], preg42_recover_table_to_gpr[9], preg41_recover_table_to_gpr[9], preg40_recover_table_to_gpr[9],
                                 preg39_recover_table_to_gpr[9], preg38_recover_table_to_gpr[9], preg37_recover_table_to_gpr[9], preg36_recover_table_to_gpr[9],
                                 preg35_recover_table_to_gpr[9], preg34_recover_table_to_gpr[9], preg33_recover_table_to_gpr[9], preg32_recover_table_to_gpr[9],
                                 preg31_recover_table_to_gpr[9], preg30_recover_table_to_gpr[9], preg29_recover_table_to_gpr[9], preg28_recover_table_to_gpr[9],
                                 preg27_recover_table_to_gpr[9], preg26_recover_table_to_gpr[9], preg25_recover_table_to_gpr[9], preg24_recover_table_to_gpr[9],
                                 preg23_recover_table_to_gpr[9], preg22_recover_table_to_gpr[9], preg21_recover_table_to_gpr[9], preg20_recover_table_to_gpr[9],
                                 preg19_recover_table_to_gpr[9], preg18_recover_table_to_gpr[9], preg17_recover_table_to_gpr[9], preg16_recover_table_to_gpr[9],
                                 preg15_recover_table_to_gpr[9], preg14_recover_table_to_gpr[9], preg13_recover_table_to_gpr[9], preg12_recover_table_to_gpr[9],
                                 preg11_recover_table_to_gpr[9], preg10_recover_table_to_gpr[9], preg9_recover_table_to_gpr[9],  preg8_recover_table_to_gpr[9] ,
                                 preg7_recover_table_to_gpr[9],  preg6_recover_table_to_gpr[9],  preg5_recover_table_to_gpr[9],  preg4_recover_table_to_gpr[9] ,
                                 preg3_recover_table_to_gpr[9],  preg2_recover_table_to_gpr[9],  preg1_recover_table_to_gpr[9],  preg0_recover_table_to_gpr[9]};
    assign gpr10_recover_table = {preg63_recover_table_to_gpr[10], preg62_recover_table_to_gpr[10], preg61_recover_table_to_gpr[10], preg60_recover_table_to_gpr[10],
                                 preg59_recover_table_to_gpr[10], preg58_recover_table_to_gpr[10], preg57_recover_table_to_gpr[10], preg56_recover_table_to_gpr[10],
                                 preg55_recover_table_to_gpr[10], preg54_recover_table_to_gpr[10], preg53_recover_table_to_gpr[10], preg52_recover_table_to_gpr[10],
                                 preg51_recover_table_to_gpr[10], preg50_recover_table_to_gpr[10], preg49_recover_table_to_gpr[10], preg48_recover_table_to_gpr[10],
                                 preg47_recover_table_to_gpr[10], preg46_recover_table_to_gpr[10], preg45_recover_table_to_gpr[10], preg44_recover_table_to_gpr[10],
                                 preg43_recover_table_to_gpr[10], preg42_recover_table_to_gpr[10], preg41_recover_table_to_gpr[10], preg40_recover_table_to_gpr[10],
                                 preg39_recover_table_to_gpr[10], preg38_recover_table_to_gpr[10], preg37_recover_table_to_gpr[10], preg36_recover_table_to_gpr[10],
                                 preg35_recover_table_to_gpr[10], preg34_recover_table_to_gpr[10], preg33_recover_table_to_gpr[10], preg32_recover_table_to_gpr[10],
                                 preg31_recover_table_to_gpr[10], preg30_recover_table_to_gpr[10], preg29_recover_table_to_gpr[10], preg28_recover_table_to_gpr[10],
                                 preg27_recover_table_to_gpr[10], preg26_recover_table_to_gpr[10], preg25_recover_table_to_gpr[10], preg24_recover_table_to_gpr[10],
                                 preg23_recover_table_to_gpr[10], preg22_recover_table_to_gpr[10], preg21_recover_table_to_gpr[10], preg20_recover_table_to_gpr[10],
                                 preg19_recover_table_to_gpr[10], preg18_recover_table_to_gpr[10], preg17_recover_table_to_gpr[10], preg16_recover_table_to_gpr[10],
                                 preg15_recover_table_to_gpr[10], preg14_recover_table_to_gpr[10], preg13_recover_table_to_gpr[10], preg12_recover_table_to_gpr[10],
                                 preg11_recover_table_to_gpr[10], preg10_recover_table_to_gpr[10], preg9_recover_table_to_gpr[10],  preg8_recover_table_to_gpr[10] ,
                                 preg7_recover_table_to_gpr[10],  preg6_recover_table_to_gpr[10],  preg5_recover_table_to_gpr[10],  preg4_recover_table_to_gpr[10] ,
                                 preg3_recover_table_to_gpr[10],  preg2_recover_table_to_gpr[10],  preg1_recover_table_to_gpr[10],  preg0_recover_table_to_gpr[10]};
    assign gpr11_recover_table = {preg63_recover_table_to_gpr[11], preg62_recover_table_to_gpr[11], preg61_recover_table_to_gpr[11], preg60_recover_table_to_gpr[11],
                                 preg59_recover_table_to_gpr[11], preg58_recover_table_to_gpr[11], preg57_recover_table_to_gpr[11], preg56_recover_table_to_gpr[11],
                                 preg55_recover_table_to_gpr[11], preg54_recover_table_to_gpr[11], preg53_recover_table_to_gpr[11], preg52_recover_table_to_gpr[11],
                                 preg51_recover_table_to_gpr[11], preg50_recover_table_to_gpr[11], preg49_recover_table_to_gpr[11], preg48_recover_table_to_gpr[11],
                                 preg47_recover_table_to_gpr[11], preg46_recover_table_to_gpr[11], preg45_recover_table_to_gpr[11], preg44_recover_table_to_gpr[11],
                                 preg43_recover_table_to_gpr[11], preg42_recover_table_to_gpr[11], preg41_recover_table_to_gpr[11], preg40_recover_table_to_gpr[11],
                                 preg39_recover_table_to_gpr[11], preg38_recover_table_to_gpr[11], preg37_recover_table_to_gpr[11], preg36_recover_table_to_gpr[11],
                                 preg35_recover_table_to_gpr[11], preg34_recover_table_to_gpr[11], preg33_recover_table_to_gpr[11], preg32_recover_table_to_gpr[11],
                                 preg31_recover_table_to_gpr[11], preg30_recover_table_to_gpr[11], preg29_recover_table_to_gpr[11], preg28_recover_table_to_gpr[11],
                                 preg27_recover_table_to_gpr[11], preg26_recover_table_to_gpr[11], preg25_recover_table_to_gpr[11], preg24_recover_table_to_gpr[11],
                                 preg23_recover_table_to_gpr[11], preg22_recover_table_to_gpr[11], preg21_recover_table_to_gpr[11], preg20_recover_table_to_gpr[11],
                                 preg19_recover_table_to_gpr[11], preg18_recover_table_to_gpr[11], preg17_recover_table_to_gpr[11], preg16_recover_table_to_gpr[11],
                                 preg15_recover_table_to_gpr[11], preg14_recover_table_to_gpr[11], preg13_recover_table_to_gpr[11], preg12_recover_table_to_gpr[11],
                                 preg11_recover_table_to_gpr[11], preg10_recover_table_to_gpr[11], preg9_recover_table_to_gpr[11],  preg8_recover_table_to_gpr[11] ,
                                 preg7_recover_table_to_gpr[11],  preg6_recover_table_to_gpr[11],  preg5_recover_table_to_gpr[11],  preg4_recover_table_to_gpr[11] ,
                                 preg3_recover_table_to_gpr[11],  preg2_recover_table_to_gpr[11],  preg1_recover_table_to_gpr[11],  preg0_recover_table_to_gpr[11]};
    assign gpr12_recover_table = {preg63_recover_table_to_gpr[12], preg62_recover_table_to_gpr[12], preg61_recover_table_to_gpr[12], preg60_recover_table_to_gpr[12],
                                 preg59_recover_table_to_gpr[12], preg58_recover_table_to_gpr[12], preg57_recover_table_to_gpr[12], preg56_recover_table_to_gpr[12],
                                 preg55_recover_table_to_gpr[12], preg54_recover_table_to_gpr[12], preg53_recover_table_to_gpr[12], preg52_recover_table_to_gpr[12],
                                 preg51_recover_table_to_gpr[12], preg50_recover_table_to_gpr[12], preg49_recover_table_to_gpr[12], preg48_recover_table_to_gpr[12],
                                 preg47_recover_table_to_gpr[12], preg46_recover_table_to_gpr[12], preg45_recover_table_to_gpr[12], preg44_recover_table_to_gpr[12],
                                 preg43_recover_table_to_gpr[12], preg42_recover_table_to_gpr[12], preg41_recover_table_to_gpr[12], preg40_recover_table_to_gpr[12],
                                 preg39_recover_table_to_gpr[12], preg38_recover_table_to_gpr[12], preg37_recover_table_to_gpr[12], preg36_recover_table_to_gpr[12],
                                 preg35_recover_table_to_gpr[12], preg34_recover_table_to_gpr[12], preg33_recover_table_to_gpr[12], preg32_recover_table_to_gpr[12],
                                 preg31_recover_table_to_gpr[12], preg30_recover_table_to_gpr[12], preg29_recover_table_to_gpr[12], preg28_recover_table_to_gpr[12],
                                 preg27_recover_table_to_gpr[12], preg26_recover_table_to_gpr[12], preg25_recover_table_to_gpr[12], preg24_recover_table_to_gpr[12],
                                 preg23_recover_table_to_gpr[12], preg22_recover_table_to_gpr[12], preg21_recover_table_to_gpr[12], preg20_recover_table_to_gpr[12],
                                 preg19_recover_table_to_gpr[12], preg18_recover_table_to_gpr[12], preg17_recover_table_to_gpr[12], preg16_recover_table_to_gpr[12],
                                 preg15_recover_table_to_gpr[12], preg14_recover_table_to_gpr[12], preg13_recover_table_to_gpr[12], preg12_recover_table_to_gpr[12],
                                 preg11_recover_table_to_gpr[12], preg10_recover_table_to_gpr[12], preg9_recover_table_to_gpr[12],  preg8_recover_table_to_gpr[12] ,
                                 preg7_recover_table_to_gpr[12],  preg6_recover_table_to_gpr[12],  preg5_recover_table_to_gpr[12],  preg4_recover_table_to_gpr[12] ,
                                 preg3_recover_table_to_gpr[12],  preg2_recover_table_to_gpr[12],  preg1_recover_table_to_gpr[12],  preg0_recover_table_to_gpr[12]};
    assign gpr13_recover_table = {preg63_recover_table_to_gpr[13], preg62_recover_table_to_gpr[13], preg61_recover_table_to_gpr[13], preg60_recover_table_to_gpr[13],
                                 preg59_recover_table_to_gpr[13], preg58_recover_table_to_gpr[13], preg57_recover_table_to_gpr[13], preg56_recover_table_to_gpr[13],
                                 preg55_recover_table_to_gpr[13], preg54_recover_table_to_gpr[13], preg53_recover_table_to_gpr[13], preg52_recover_table_to_gpr[13],
                                 preg51_recover_table_to_gpr[13], preg50_recover_table_to_gpr[13], preg49_recover_table_to_gpr[13], preg48_recover_table_to_gpr[13],
                                 preg47_recover_table_to_gpr[13], preg46_recover_table_to_gpr[13], preg45_recover_table_to_gpr[13], preg44_recover_table_to_gpr[13],
                                 preg43_recover_table_to_gpr[13], preg42_recover_table_to_gpr[13], preg41_recover_table_to_gpr[13], preg40_recover_table_to_gpr[13],
                                 preg39_recover_table_to_gpr[13], preg38_recover_table_to_gpr[13], preg37_recover_table_to_gpr[13], preg36_recover_table_to_gpr[13],
                                 preg35_recover_table_to_gpr[13], preg34_recover_table_to_gpr[13], preg33_recover_table_to_gpr[13], preg32_recover_table_to_gpr[13],
                                 preg31_recover_table_to_gpr[13], preg30_recover_table_to_gpr[13], preg29_recover_table_to_gpr[13], preg28_recover_table_to_gpr[13],
                                 preg27_recover_table_to_gpr[13], preg26_recover_table_to_gpr[13], preg25_recover_table_to_gpr[13], preg24_recover_table_to_gpr[13],
                                 preg23_recover_table_to_gpr[13], preg22_recover_table_to_gpr[13], preg21_recover_table_to_gpr[13], preg20_recover_table_to_gpr[13],
                                 preg19_recover_table_to_gpr[13], preg18_recover_table_to_gpr[13], preg17_recover_table_to_gpr[13], preg16_recover_table_to_gpr[13],
                                 preg15_recover_table_to_gpr[13], preg14_recover_table_to_gpr[13], preg13_recover_table_to_gpr[13], preg12_recover_table_to_gpr[13],
                                 preg11_recover_table_to_gpr[13], preg10_recover_table_to_gpr[13], preg9_recover_table_to_gpr[13],  preg8_recover_table_to_gpr[13] ,
                                 preg7_recover_table_to_gpr[13],  preg6_recover_table_to_gpr[13],  preg5_recover_table_to_gpr[13],  preg4_recover_table_to_gpr[13] ,
                                 preg3_recover_table_to_gpr[13],  preg2_recover_table_to_gpr[13],  preg1_recover_table_to_gpr[13],  preg0_recover_table_to_gpr[13]};
    assign gpr14_recover_table = {preg63_recover_table_to_gpr[14], preg62_recover_table_to_gpr[14], preg61_recover_table_to_gpr[14], preg60_recover_table_to_gpr[14],
                                 preg59_recover_table_to_gpr[14], preg58_recover_table_to_gpr[14], preg57_recover_table_to_gpr[14], preg56_recover_table_to_gpr[14],
                                 preg55_recover_table_to_gpr[14], preg54_recover_table_to_gpr[14], preg53_recover_table_to_gpr[14], preg52_recover_table_to_gpr[14],
                                 preg51_recover_table_to_gpr[14], preg50_recover_table_to_gpr[14], preg49_recover_table_to_gpr[14], preg48_recover_table_to_gpr[14],
                                 preg47_recover_table_to_gpr[14], preg46_recover_table_to_gpr[14], preg45_recover_table_to_gpr[14], preg44_recover_table_to_gpr[14],
                                 preg43_recover_table_to_gpr[14], preg42_recover_table_to_gpr[14], preg41_recover_table_to_gpr[14], preg40_recover_table_to_gpr[14],
                                 preg39_recover_table_to_gpr[14], preg38_recover_table_to_gpr[14], preg37_recover_table_to_gpr[14], preg36_recover_table_to_gpr[14],
                                 preg35_recover_table_to_gpr[14], preg34_recover_table_to_gpr[14], preg33_recover_table_to_gpr[14], preg32_recover_table_to_gpr[14],
                                 preg31_recover_table_to_gpr[14], preg30_recover_table_to_gpr[14], preg29_recover_table_to_gpr[14], preg28_recover_table_to_gpr[14],
                                 preg27_recover_table_to_gpr[14], preg26_recover_table_to_gpr[14], preg25_recover_table_to_gpr[14], preg24_recover_table_to_gpr[14],
                                 preg23_recover_table_to_gpr[14], preg22_recover_table_to_gpr[14], preg21_recover_table_to_gpr[14], preg20_recover_table_to_gpr[14],
                                 preg19_recover_table_to_gpr[14], preg18_recover_table_to_gpr[14], preg17_recover_table_to_gpr[14], preg16_recover_table_to_gpr[14],
                                 preg15_recover_table_to_gpr[14], preg14_recover_table_to_gpr[14], preg13_recover_table_to_gpr[14], preg12_recover_table_to_gpr[14],
                                 preg11_recover_table_to_gpr[14], preg10_recover_table_to_gpr[14], preg9_recover_table_to_gpr[14],  preg8_recover_table_to_gpr[14] ,
                                 preg7_recover_table_to_gpr[14],  preg6_recover_table_to_gpr[14],  preg5_recover_table_to_gpr[14],  preg4_recover_table_to_gpr[14] ,
                                 preg3_recover_table_to_gpr[14],  preg2_recover_table_to_gpr[14],  preg1_recover_table_to_gpr[14],  preg0_recover_table_to_gpr[14]};
    assign gpr15_recover_table = {preg63_recover_table_to_gpr[15], preg62_recover_table_to_gpr[15], preg61_recover_table_to_gpr[15], preg60_recover_table_to_gpr[15],
                                 preg59_recover_table_to_gpr[15], preg58_recover_table_to_gpr[15], preg57_recover_table_to_gpr[15], preg56_recover_table_to_gpr[15],
                                 preg55_recover_table_to_gpr[15], preg54_recover_table_to_gpr[15], preg53_recover_table_to_gpr[15], preg52_recover_table_to_gpr[15],
                                 preg51_recover_table_to_gpr[15], preg50_recover_table_to_gpr[15], preg49_recover_table_to_gpr[15], preg48_recover_table_to_gpr[15],
                                 preg47_recover_table_to_gpr[15], preg46_recover_table_to_gpr[15], preg45_recover_table_to_gpr[15], preg44_recover_table_to_gpr[15],
                                 preg43_recover_table_to_gpr[15], preg42_recover_table_to_gpr[15], preg41_recover_table_to_gpr[15], preg40_recover_table_to_gpr[15],
                                 preg39_recover_table_to_gpr[15], preg38_recover_table_to_gpr[15], preg37_recover_table_to_gpr[15], preg36_recover_table_to_gpr[15],
                                 preg35_recover_table_to_gpr[15], preg34_recover_table_to_gpr[15], preg33_recover_table_to_gpr[15], preg32_recover_table_to_gpr[15],
                                 preg31_recover_table_to_gpr[15], preg30_recover_table_to_gpr[15], preg29_recover_table_to_gpr[15], preg28_recover_table_to_gpr[15],
                                 preg27_recover_table_to_gpr[15], preg26_recover_table_to_gpr[15], preg25_recover_table_to_gpr[15], preg24_recover_table_to_gpr[15],
                                 preg23_recover_table_to_gpr[15], preg22_recover_table_to_gpr[15], preg21_recover_table_to_gpr[15], preg20_recover_table_to_gpr[15],
                                 preg19_recover_table_to_gpr[15], preg18_recover_table_to_gpr[15], preg17_recover_table_to_gpr[15], preg16_recover_table_to_gpr[15],
                                 preg15_recover_table_to_gpr[15], preg14_recover_table_to_gpr[15], preg13_recover_table_to_gpr[15], preg12_recover_table_to_gpr[15],
                                 preg11_recover_table_to_gpr[15], preg10_recover_table_to_gpr[15], preg9_recover_table_to_gpr[15],  preg8_recover_table_to_gpr[15] ,
                                 preg7_recover_table_to_gpr[15],  preg6_recover_table_to_gpr[15],  preg5_recover_table_to_gpr[15],  preg4_recover_table_to_gpr[15] ,
                                 preg3_recover_table_to_gpr[15],  preg2_recover_table_to_gpr[15],  preg1_recover_table_to_gpr[15],  preg0_recover_table_to_gpr[15]};
    assign gpr16_recover_table = {preg63_recover_table_to_gpr[16], preg62_recover_table_to_gpr[16], preg61_recover_table_to_gpr[16], preg60_recover_table_to_gpr[16],
                                 preg59_recover_table_to_gpr[16], preg58_recover_table_to_gpr[16], preg57_recover_table_to_gpr[16], preg56_recover_table_to_gpr[16],
                                 preg55_recover_table_to_gpr[16], preg54_recover_table_to_gpr[16], preg53_recover_table_to_gpr[16], preg52_recover_table_to_gpr[16],
                                 preg51_recover_table_to_gpr[16], preg50_recover_table_to_gpr[16], preg49_recover_table_to_gpr[16], preg48_recover_table_to_gpr[16],
                                 preg47_recover_table_to_gpr[16], preg46_recover_table_to_gpr[16], preg45_recover_table_to_gpr[16], preg44_recover_table_to_gpr[16],
                                 preg43_recover_table_to_gpr[16], preg42_recover_table_to_gpr[16], preg41_recover_table_to_gpr[16], preg40_recover_table_to_gpr[16],
                                 preg39_recover_table_to_gpr[16], preg38_recover_table_to_gpr[16], preg37_recover_table_to_gpr[16], preg36_recover_table_to_gpr[16],
                                 preg35_recover_table_to_gpr[16], preg34_recover_table_to_gpr[16], preg33_recover_table_to_gpr[16], preg32_recover_table_to_gpr[16],
                                 preg31_recover_table_to_gpr[16], preg30_recover_table_to_gpr[16], preg29_recover_table_to_gpr[16], preg28_recover_table_to_gpr[16],
                                 preg27_recover_table_to_gpr[16], preg26_recover_table_to_gpr[16], preg25_recover_table_to_gpr[16], preg24_recover_table_to_gpr[16],
                                 preg23_recover_table_to_gpr[16], preg22_recover_table_to_gpr[16], preg21_recover_table_to_gpr[16], preg20_recover_table_to_gpr[16],
                                 preg19_recover_table_to_gpr[16], preg18_recover_table_to_gpr[16], preg17_recover_table_to_gpr[16], preg16_recover_table_to_gpr[16],
                                 preg15_recover_table_to_gpr[16], preg14_recover_table_to_gpr[16], preg13_recover_table_to_gpr[16], preg12_recover_table_to_gpr[16],
                                 preg11_recover_table_to_gpr[16], preg10_recover_table_to_gpr[16], preg9_recover_table_to_gpr[16],  preg8_recover_table_to_gpr[16] ,
                                 preg7_recover_table_to_gpr[16],  preg6_recover_table_to_gpr[16],  preg5_recover_table_to_gpr[16],  preg4_recover_table_to_gpr[16] ,
                                 preg3_recover_table_to_gpr[16],  preg2_recover_table_to_gpr[16],  preg1_recover_table_to_gpr[16],  preg0_recover_table_to_gpr[16]};
    assign gpr17_recover_table = {preg63_recover_table_to_gpr[17], preg62_recover_table_to_gpr[17], preg61_recover_table_to_gpr[17], preg60_recover_table_to_gpr[17],
                                 preg59_recover_table_to_gpr[17], preg58_recover_table_to_gpr[17], preg57_recover_table_to_gpr[17], preg56_recover_table_to_gpr[17],
                                 preg55_recover_table_to_gpr[17], preg54_recover_table_to_gpr[17], preg53_recover_table_to_gpr[17], preg52_recover_table_to_gpr[17],
                                 preg51_recover_table_to_gpr[17], preg50_recover_table_to_gpr[17], preg49_recover_table_to_gpr[17], preg48_recover_table_to_gpr[17],
                                 preg47_recover_table_to_gpr[17], preg46_recover_table_to_gpr[17], preg45_recover_table_to_gpr[17], preg44_recover_table_to_gpr[17],
                                 preg43_recover_table_to_gpr[17], preg42_recover_table_to_gpr[17], preg41_recover_table_to_gpr[17], preg40_recover_table_to_gpr[17],
                                 preg39_recover_table_to_gpr[17], preg38_recover_table_to_gpr[17], preg37_recover_table_to_gpr[17], preg36_recover_table_to_gpr[17],
                                 preg35_recover_table_to_gpr[17], preg34_recover_table_to_gpr[17], preg33_recover_table_to_gpr[17], preg32_recover_table_to_gpr[17],
                                 preg31_recover_table_to_gpr[17], preg30_recover_table_to_gpr[17], preg29_recover_table_to_gpr[17], preg28_recover_table_to_gpr[17],
                                 preg27_recover_table_to_gpr[17], preg26_recover_table_to_gpr[17], preg25_recover_table_to_gpr[17], preg24_recover_table_to_gpr[17],
                                 preg23_recover_table_to_gpr[17], preg22_recover_table_to_gpr[17], preg21_recover_table_to_gpr[17], preg20_recover_table_to_gpr[17],
                                 preg19_recover_table_to_gpr[17], preg18_recover_table_to_gpr[17], preg17_recover_table_to_gpr[17], preg16_recover_table_to_gpr[17],
                                 preg15_recover_table_to_gpr[17], preg14_recover_table_to_gpr[17], preg13_recover_table_to_gpr[17], preg12_recover_table_to_gpr[17],
                                 preg11_recover_table_to_gpr[17], preg10_recover_table_to_gpr[17], preg9_recover_table_to_gpr[17],  preg8_recover_table_to_gpr[17] ,
                                 preg7_recover_table_to_gpr[17],  preg6_recover_table_to_gpr[17],  preg5_recover_table_to_gpr[17],  preg4_recover_table_to_gpr[17] ,
                                 preg3_recover_table_to_gpr[17],  preg2_recover_table_to_gpr[17],  preg1_recover_table_to_gpr[17],  preg0_recover_table_to_gpr[17]};
    assign gpr18_recover_table = {preg63_recover_table_to_gpr[18], preg62_recover_table_to_gpr[18], preg61_recover_table_to_gpr[18], preg60_recover_table_to_gpr[18],
                                 preg59_recover_table_to_gpr[18], preg58_recover_table_to_gpr[18], preg57_recover_table_to_gpr[18], preg56_recover_table_to_gpr[18],
                                 preg55_recover_table_to_gpr[18], preg54_recover_table_to_gpr[18], preg53_recover_table_to_gpr[18], preg52_recover_table_to_gpr[18],
                                 preg51_recover_table_to_gpr[18], preg50_recover_table_to_gpr[18], preg49_recover_table_to_gpr[18], preg48_recover_table_to_gpr[18],
                                 preg47_recover_table_to_gpr[18], preg46_recover_table_to_gpr[18], preg45_recover_table_to_gpr[18], preg44_recover_table_to_gpr[18],
                                 preg43_recover_table_to_gpr[18], preg42_recover_table_to_gpr[18], preg41_recover_table_to_gpr[18], preg40_recover_table_to_gpr[18],
                                 preg39_recover_table_to_gpr[18], preg38_recover_table_to_gpr[18], preg37_recover_table_to_gpr[18], preg36_recover_table_to_gpr[18],
                                 preg35_recover_table_to_gpr[18], preg34_recover_table_to_gpr[18], preg33_recover_table_to_gpr[18], preg32_recover_table_to_gpr[18],
                                 preg31_recover_table_to_gpr[18], preg30_recover_table_to_gpr[18], preg29_recover_table_to_gpr[18], preg28_recover_table_to_gpr[18],
                                 preg27_recover_table_to_gpr[18], preg26_recover_table_to_gpr[18], preg25_recover_table_to_gpr[18], preg24_recover_table_to_gpr[18],
                                 preg23_recover_table_to_gpr[18], preg22_recover_table_to_gpr[18], preg21_recover_table_to_gpr[18], preg20_recover_table_to_gpr[18],
                                 preg19_recover_table_to_gpr[18], preg18_recover_table_to_gpr[18], preg17_recover_table_to_gpr[18], preg16_recover_table_to_gpr[18],
                                 preg15_recover_table_to_gpr[18], preg14_recover_table_to_gpr[18], preg13_recover_table_to_gpr[18], preg12_recover_table_to_gpr[18],
                                 preg11_recover_table_to_gpr[18], preg10_recover_table_to_gpr[18], preg9_recover_table_to_gpr[18],  preg8_recover_table_to_gpr[18] ,
                                 preg7_recover_table_to_gpr[18],  preg6_recover_table_to_gpr[18],  preg5_recover_table_to_gpr[18],  preg4_recover_table_to_gpr[18] ,
                                 preg3_recover_table_to_gpr[18],  preg2_recover_table_to_gpr[18],  preg1_recover_table_to_gpr[18],  preg0_recover_table_to_gpr[18]};
    assign gpr19_recover_table = {preg63_recover_table_to_gpr[19], preg62_recover_table_to_gpr[19], preg61_recover_table_to_gpr[19], preg60_recover_table_to_gpr[19],
                                 preg59_recover_table_to_gpr[19], preg58_recover_table_to_gpr[19], preg57_recover_table_to_gpr[19], preg56_recover_table_to_gpr[19],
                                 preg55_recover_table_to_gpr[19], preg54_recover_table_to_gpr[19], preg53_recover_table_to_gpr[19], preg52_recover_table_to_gpr[19],
                                 preg51_recover_table_to_gpr[19], preg50_recover_table_to_gpr[19], preg49_recover_table_to_gpr[19], preg48_recover_table_to_gpr[19],
                                 preg47_recover_table_to_gpr[19], preg46_recover_table_to_gpr[19], preg45_recover_table_to_gpr[19], preg44_recover_table_to_gpr[19],
                                 preg43_recover_table_to_gpr[19], preg42_recover_table_to_gpr[19], preg41_recover_table_to_gpr[19], preg40_recover_table_to_gpr[19],
                                 preg39_recover_table_to_gpr[19], preg38_recover_table_to_gpr[19], preg37_recover_table_to_gpr[19], preg36_recover_table_to_gpr[19],
                                 preg35_recover_table_to_gpr[19], preg34_recover_table_to_gpr[19], preg33_recover_table_to_gpr[19], preg32_recover_table_to_gpr[19],
                                 preg31_recover_table_to_gpr[19], preg30_recover_table_to_gpr[19], preg29_recover_table_to_gpr[19], preg28_recover_table_to_gpr[19],
                                 preg27_recover_table_to_gpr[19], preg26_recover_table_to_gpr[19], preg25_recover_table_to_gpr[19], preg24_recover_table_to_gpr[19],
                                 preg23_recover_table_to_gpr[19], preg22_recover_table_to_gpr[19], preg21_recover_table_to_gpr[19], preg20_recover_table_to_gpr[19],
                                 preg19_recover_table_to_gpr[19], preg18_recover_table_to_gpr[19], preg17_recover_table_to_gpr[19], preg16_recover_table_to_gpr[19],
                                 preg15_recover_table_to_gpr[19], preg14_recover_table_to_gpr[19], preg13_recover_table_to_gpr[19], preg12_recover_table_to_gpr[19],
                                 preg11_recover_table_to_gpr[19], preg10_recover_table_to_gpr[19], preg9_recover_table_to_gpr[19],  preg8_recover_table_to_gpr[19] ,
                                 preg7_recover_table_to_gpr[19],  preg6_recover_table_to_gpr[19],  preg5_recover_table_to_gpr[19],  preg4_recover_table_to_gpr[19] ,
                                 preg3_recover_table_to_gpr[19],  preg2_recover_table_to_gpr[19],  preg1_recover_table_to_gpr[19],  preg0_recover_table_to_gpr[19]};
    assign gpr20_recover_table = {preg63_recover_table_to_gpr[20], preg62_recover_table_to_gpr[20], preg61_recover_table_to_gpr[20], preg60_recover_table_to_gpr[20],
                                 preg59_recover_table_to_gpr[20], preg58_recover_table_to_gpr[20], preg57_recover_table_to_gpr[20], preg56_recover_table_to_gpr[20],
                                 preg55_recover_table_to_gpr[20], preg54_recover_table_to_gpr[20], preg53_recover_table_to_gpr[20], preg52_recover_table_to_gpr[20],
                                 preg51_recover_table_to_gpr[20], preg50_recover_table_to_gpr[20], preg49_recover_table_to_gpr[20], preg48_recover_table_to_gpr[20],
                                 preg47_recover_table_to_gpr[20], preg46_recover_table_to_gpr[20], preg45_recover_table_to_gpr[20], preg44_recover_table_to_gpr[20],
                                 preg43_recover_table_to_gpr[20], preg42_recover_table_to_gpr[20], preg41_recover_table_to_gpr[20], preg40_recover_table_to_gpr[20],
                                 preg39_recover_table_to_gpr[20], preg38_recover_table_to_gpr[20], preg37_recover_table_to_gpr[20], preg36_recover_table_to_gpr[20],
                                 preg35_recover_table_to_gpr[20], preg34_recover_table_to_gpr[20], preg33_recover_table_to_gpr[20], preg32_recover_table_to_gpr[20],
                                 preg31_recover_table_to_gpr[20], preg30_recover_table_to_gpr[20], preg29_recover_table_to_gpr[20], preg28_recover_table_to_gpr[20],
                                 preg27_recover_table_to_gpr[20], preg26_recover_table_to_gpr[20], preg25_recover_table_to_gpr[20], preg24_recover_table_to_gpr[20],
                                 preg23_recover_table_to_gpr[20], preg22_recover_table_to_gpr[20], preg21_recover_table_to_gpr[20], preg20_recover_table_to_gpr[20],
                                 preg19_recover_table_to_gpr[20], preg18_recover_table_to_gpr[20], preg17_recover_table_to_gpr[20], preg16_recover_table_to_gpr[20],
                                 preg15_recover_table_to_gpr[20], preg14_recover_table_to_gpr[20], preg13_recover_table_to_gpr[20], preg12_recover_table_to_gpr[20],
                                 preg11_recover_table_to_gpr[20], preg10_recover_table_to_gpr[20], preg9_recover_table_to_gpr[20],  preg8_recover_table_to_gpr[20] ,
                                 preg7_recover_table_to_gpr[20],  preg6_recover_table_to_gpr[20],  preg5_recover_table_to_gpr[20],  preg4_recover_table_to_gpr[20] ,
                                 preg3_recover_table_to_gpr[20],  preg2_recover_table_to_gpr[20],  preg1_recover_table_to_gpr[20],  preg0_recover_table_to_gpr[20]};
    assign gpr21_recover_table = {preg63_recover_table_to_gpr[21], preg62_recover_table_to_gpr[21], preg61_recover_table_to_gpr[21], preg60_recover_table_to_gpr[21],
                                 preg59_recover_table_to_gpr[21], preg58_recover_table_to_gpr[21], preg57_recover_table_to_gpr[21], preg56_recover_table_to_gpr[21],
                                 preg55_recover_table_to_gpr[21], preg54_recover_table_to_gpr[21], preg53_recover_table_to_gpr[21], preg52_recover_table_to_gpr[21],
                                 preg51_recover_table_to_gpr[21], preg50_recover_table_to_gpr[21], preg49_recover_table_to_gpr[21], preg48_recover_table_to_gpr[21],
                                 preg47_recover_table_to_gpr[21], preg46_recover_table_to_gpr[21], preg45_recover_table_to_gpr[21], preg44_recover_table_to_gpr[21],
                                 preg43_recover_table_to_gpr[21], preg42_recover_table_to_gpr[21], preg41_recover_table_to_gpr[21], preg40_recover_table_to_gpr[21],
                                 preg39_recover_table_to_gpr[21], preg38_recover_table_to_gpr[21], preg37_recover_table_to_gpr[21], preg36_recover_table_to_gpr[21],
                                 preg35_recover_table_to_gpr[21], preg34_recover_table_to_gpr[21], preg33_recover_table_to_gpr[21], preg32_recover_table_to_gpr[21],
                                 preg31_recover_table_to_gpr[21], preg30_recover_table_to_gpr[21], preg29_recover_table_to_gpr[21], preg28_recover_table_to_gpr[21],
                                 preg27_recover_table_to_gpr[21], preg26_recover_table_to_gpr[21], preg25_recover_table_to_gpr[21], preg24_recover_table_to_gpr[21],
                                 preg23_recover_table_to_gpr[21], preg22_recover_table_to_gpr[21], preg21_recover_table_to_gpr[21], preg20_recover_table_to_gpr[21],
                                 preg19_recover_table_to_gpr[21], preg18_recover_table_to_gpr[21], preg17_recover_table_to_gpr[21], preg16_recover_table_to_gpr[21],
                                 preg15_recover_table_to_gpr[21], preg14_recover_table_to_gpr[21], preg13_recover_table_to_gpr[21], preg12_recover_table_to_gpr[21],
                                 preg11_recover_table_to_gpr[21], preg10_recover_table_to_gpr[21], preg9_recover_table_to_gpr[21],  preg8_recover_table_to_gpr[21] ,
                                 preg7_recover_table_to_gpr[21],  preg6_recover_table_to_gpr[21],  preg5_recover_table_to_gpr[21],  preg4_recover_table_to_gpr[21] ,
                                 preg3_recover_table_to_gpr[21],  preg2_recover_table_to_gpr[21],  preg1_recover_table_to_gpr[21],  preg0_recover_table_to_gpr[21]};
    assign gpr22_recover_table = {preg63_recover_table_to_gpr[22], preg62_recover_table_to_gpr[22], preg61_recover_table_to_gpr[22], preg60_recover_table_to_gpr[22],
                                 preg59_recover_table_to_gpr[22], preg58_recover_table_to_gpr[22], preg57_recover_table_to_gpr[22], preg56_recover_table_to_gpr[22],
                                 preg55_recover_table_to_gpr[22], preg54_recover_table_to_gpr[22], preg53_recover_table_to_gpr[22], preg52_recover_table_to_gpr[22],
                                 preg51_recover_table_to_gpr[22], preg50_recover_table_to_gpr[22], preg49_recover_table_to_gpr[22], preg48_recover_table_to_gpr[22],
                                 preg47_recover_table_to_gpr[22], preg46_recover_table_to_gpr[22], preg45_recover_table_to_gpr[22], preg44_recover_table_to_gpr[22],
                                 preg43_recover_table_to_gpr[22], preg42_recover_table_to_gpr[22], preg41_recover_table_to_gpr[22], preg40_recover_table_to_gpr[22],
                                 preg39_recover_table_to_gpr[22], preg38_recover_table_to_gpr[22], preg37_recover_table_to_gpr[22], preg36_recover_table_to_gpr[22],
                                 preg35_recover_table_to_gpr[22], preg34_recover_table_to_gpr[22], preg33_recover_table_to_gpr[22], preg32_recover_table_to_gpr[22],
                                 preg31_recover_table_to_gpr[22], preg30_recover_table_to_gpr[22], preg29_recover_table_to_gpr[22], preg28_recover_table_to_gpr[22],
                                 preg27_recover_table_to_gpr[22], preg26_recover_table_to_gpr[22], preg25_recover_table_to_gpr[22], preg24_recover_table_to_gpr[22],
                                 preg23_recover_table_to_gpr[22], preg22_recover_table_to_gpr[22], preg21_recover_table_to_gpr[22], preg20_recover_table_to_gpr[22],
                                 preg19_recover_table_to_gpr[22], preg18_recover_table_to_gpr[22], preg17_recover_table_to_gpr[22], preg16_recover_table_to_gpr[22],
                                 preg15_recover_table_to_gpr[22], preg14_recover_table_to_gpr[22], preg13_recover_table_to_gpr[22], preg12_recover_table_to_gpr[22],
                                 preg11_recover_table_to_gpr[22], preg10_recover_table_to_gpr[22], preg9_recover_table_to_gpr[22],  preg8_recover_table_to_gpr[22] ,
                                 preg7_recover_table_to_gpr[22],  preg6_recover_table_to_gpr[22],  preg5_recover_table_to_gpr[22],  preg4_recover_table_to_gpr[22] ,
                                 preg3_recover_table_to_gpr[22],  preg2_recover_table_to_gpr[22],  preg1_recover_table_to_gpr[22],  preg0_recover_table_to_gpr[22]};
    assign gpr23_recover_table = {preg63_recover_table_to_gpr[23], preg62_recover_table_to_gpr[23], preg61_recover_table_to_gpr[23], preg60_recover_table_to_gpr[23],
                                 preg59_recover_table_to_gpr[23], preg58_recover_table_to_gpr[23], preg57_recover_table_to_gpr[23], preg56_recover_table_to_gpr[23],
                                 preg55_recover_table_to_gpr[23], preg54_recover_table_to_gpr[23], preg53_recover_table_to_gpr[23], preg52_recover_table_to_gpr[23],
                                 preg51_recover_table_to_gpr[23], preg50_recover_table_to_gpr[23], preg49_recover_table_to_gpr[23], preg48_recover_table_to_gpr[23],
                                 preg47_recover_table_to_gpr[23], preg46_recover_table_to_gpr[23], preg45_recover_table_to_gpr[23], preg44_recover_table_to_gpr[23],
                                 preg43_recover_table_to_gpr[23], preg42_recover_table_to_gpr[23], preg41_recover_table_to_gpr[23], preg40_recover_table_to_gpr[23],
                                 preg39_recover_table_to_gpr[23], preg38_recover_table_to_gpr[23], preg37_recover_table_to_gpr[23], preg36_recover_table_to_gpr[23],
                                 preg35_recover_table_to_gpr[23], preg34_recover_table_to_gpr[23], preg33_recover_table_to_gpr[23], preg32_recover_table_to_gpr[23],
                                 preg31_recover_table_to_gpr[23], preg30_recover_table_to_gpr[23], preg29_recover_table_to_gpr[23], preg28_recover_table_to_gpr[23],
                                 preg27_recover_table_to_gpr[23], preg26_recover_table_to_gpr[23], preg25_recover_table_to_gpr[23], preg24_recover_table_to_gpr[23],
                                 preg23_recover_table_to_gpr[23], preg22_recover_table_to_gpr[23], preg21_recover_table_to_gpr[23], preg20_recover_table_to_gpr[23],
                                 preg19_recover_table_to_gpr[23], preg18_recover_table_to_gpr[23], preg17_recover_table_to_gpr[23], preg16_recover_table_to_gpr[23],
                                 preg15_recover_table_to_gpr[23], preg14_recover_table_to_gpr[23], preg13_recover_table_to_gpr[23], preg12_recover_table_to_gpr[23],
                                 preg11_recover_table_to_gpr[23], preg10_recover_table_to_gpr[23], preg9_recover_table_to_gpr[23],  preg8_recover_table_to_gpr[23] ,
                                 preg7_recover_table_to_gpr[23],  preg6_recover_table_to_gpr[23],  preg5_recover_table_to_gpr[23],  preg4_recover_table_to_gpr[23] ,
                                 preg3_recover_table_to_gpr[23],  preg2_recover_table_to_gpr[23],  preg1_recover_table_to_gpr[23],  preg0_recover_table_to_gpr[23]};
    assign gpr24_recover_table = {preg63_recover_table_to_gpr[24], preg62_recover_table_to_gpr[24], preg61_recover_table_to_gpr[24], preg60_recover_table_to_gpr[24],
                                 preg59_recover_table_to_gpr[24], preg58_recover_table_to_gpr[24], preg57_recover_table_to_gpr[24], preg56_recover_table_to_gpr[24],
                                 preg55_recover_table_to_gpr[24], preg54_recover_table_to_gpr[24], preg53_recover_table_to_gpr[24], preg52_recover_table_to_gpr[24],
                                 preg51_recover_table_to_gpr[24], preg50_recover_table_to_gpr[24], preg49_recover_table_to_gpr[24], preg48_recover_table_to_gpr[24],
                                 preg47_recover_table_to_gpr[24], preg46_recover_table_to_gpr[24], preg45_recover_table_to_gpr[24], preg44_recover_table_to_gpr[24],
                                 preg43_recover_table_to_gpr[24], preg42_recover_table_to_gpr[24], preg41_recover_table_to_gpr[24], preg40_recover_table_to_gpr[24],
                                 preg39_recover_table_to_gpr[24], preg38_recover_table_to_gpr[24], preg37_recover_table_to_gpr[24], preg36_recover_table_to_gpr[24],
                                 preg35_recover_table_to_gpr[24], preg34_recover_table_to_gpr[24], preg33_recover_table_to_gpr[24], preg32_recover_table_to_gpr[24],
                                 preg31_recover_table_to_gpr[24], preg30_recover_table_to_gpr[24], preg29_recover_table_to_gpr[24], preg28_recover_table_to_gpr[24],
                                 preg27_recover_table_to_gpr[24], preg26_recover_table_to_gpr[24], preg25_recover_table_to_gpr[24], preg24_recover_table_to_gpr[24],
                                 preg23_recover_table_to_gpr[24], preg22_recover_table_to_gpr[24], preg21_recover_table_to_gpr[24], preg20_recover_table_to_gpr[24],
                                 preg19_recover_table_to_gpr[24], preg18_recover_table_to_gpr[24], preg17_recover_table_to_gpr[24], preg16_recover_table_to_gpr[24],
                                 preg15_recover_table_to_gpr[24], preg14_recover_table_to_gpr[24], preg13_recover_table_to_gpr[24], preg12_recover_table_to_gpr[24],
                                 preg11_recover_table_to_gpr[24], preg10_recover_table_to_gpr[24], preg9_recover_table_to_gpr[24],  preg8_recover_table_to_gpr[24] ,
                                 preg7_recover_table_to_gpr[24],  preg6_recover_table_to_gpr[24],  preg5_recover_table_to_gpr[24],  preg4_recover_table_to_gpr[24] ,
                                 preg3_recover_table_to_gpr[24],  preg2_recover_table_to_gpr[24],  preg1_recover_table_to_gpr[24],  preg0_recover_table_to_gpr[24]};
    assign gpr25_recover_table = {preg63_recover_table_to_gpr[25], preg62_recover_table_to_gpr[25], preg61_recover_table_to_gpr[25], preg60_recover_table_to_gpr[25],
                                 preg59_recover_table_to_gpr[25], preg58_recover_table_to_gpr[25], preg57_recover_table_to_gpr[25], preg56_recover_table_to_gpr[25],
                                 preg55_recover_table_to_gpr[25], preg54_recover_table_to_gpr[25], preg53_recover_table_to_gpr[25], preg52_recover_table_to_gpr[25],
                                 preg51_recover_table_to_gpr[25], preg50_recover_table_to_gpr[25], preg49_recover_table_to_gpr[25], preg48_recover_table_to_gpr[25],
                                 preg47_recover_table_to_gpr[25], preg46_recover_table_to_gpr[25], preg45_recover_table_to_gpr[25], preg44_recover_table_to_gpr[25],
                                 preg43_recover_table_to_gpr[25], preg42_recover_table_to_gpr[25], preg41_recover_table_to_gpr[25], preg40_recover_table_to_gpr[25],
                                 preg39_recover_table_to_gpr[25], preg38_recover_table_to_gpr[25], preg37_recover_table_to_gpr[25], preg36_recover_table_to_gpr[25],
                                 preg35_recover_table_to_gpr[25], preg34_recover_table_to_gpr[25], preg33_recover_table_to_gpr[25], preg32_recover_table_to_gpr[25],
                                 preg31_recover_table_to_gpr[25], preg30_recover_table_to_gpr[25], preg29_recover_table_to_gpr[25], preg28_recover_table_to_gpr[25],
                                 preg27_recover_table_to_gpr[25], preg26_recover_table_to_gpr[25], preg25_recover_table_to_gpr[25], preg24_recover_table_to_gpr[25],
                                 preg23_recover_table_to_gpr[25], preg22_recover_table_to_gpr[25], preg21_recover_table_to_gpr[25], preg20_recover_table_to_gpr[25],
                                 preg19_recover_table_to_gpr[25], preg18_recover_table_to_gpr[25], preg17_recover_table_to_gpr[25], preg16_recover_table_to_gpr[25],
                                 preg15_recover_table_to_gpr[25], preg14_recover_table_to_gpr[25], preg13_recover_table_to_gpr[25], preg12_recover_table_to_gpr[25],
                                 preg11_recover_table_to_gpr[25], preg10_recover_table_to_gpr[25], preg9_recover_table_to_gpr[25],  preg8_recover_table_to_gpr[25] ,
                                 preg7_recover_table_to_gpr[25],  preg6_recover_table_to_gpr[25],  preg5_recover_table_to_gpr[25],  preg4_recover_table_to_gpr[25] ,
                                 preg3_recover_table_to_gpr[25],  preg2_recover_table_to_gpr[25],  preg1_recover_table_to_gpr[25],  preg0_recover_table_to_gpr[25]};
    assign gpr26_recover_table = {preg63_recover_table_to_gpr[26], preg62_recover_table_to_gpr[26], preg61_recover_table_to_gpr[26], preg60_recover_table_to_gpr[26],
                                 preg59_recover_table_to_gpr[26], preg58_recover_table_to_gpr[26], preg57_recover_table_to_gpr[26], preg56_recover_table_to_gpr[26],
                                 preg55_recover_table_to_gpr[26], preg54_recover_table_to_gpr[26], preg53_recover_table_to_gpr[26], preg52_recover_table_to_gpr[26],
                                 preg51_recover_table_to_gpr[26], preg50_recover_table_to_gpr[26], preg49_recover_table_to_gpr[26], preg48_recover_table_to_gpr[26],
                                 preg47_recover_table_to_gpr[26], preg46_recover_table_to_gpr[26], preg45_recover_table_to_gpr[26], preg44_recover_table_to_gpr[26],
                                 preg43_recover_table_to_gpr[26], preg42_recover_table_to_gpr[26], preg41_recover_table_to_gpr[26], preg40_recover_table_to_gpr[26],
                                 preg39_recover_table_to_gpr[26], preg38_recover_table_to_gpr[26], preg37_recover_table_to_gpr[26], preg36_recover_table_to_gpr[26],
                                 preg35_recover_table_to_gpr[26], preg34_recover_table_to_gpr[26], preg33_recover_table_to_gpr[26], preg32_recover_table_to_gpr[26],
                                 preg31_recover_table_to_gpr[26], preg30_recover_table_to_gpr[26], preg29_recover_table_to_gpr[26], preg28_recover_table_to_gpr[26],
                                 preg27_recover_table_to_gpr[26], preg26_recover_table_to_gpr[26], preg25_recover_table_to_gpr[26], preg24_recover_table_to_gpr[26],
                                 preg23_recover_table_to_gpr[26], preg22_recover_table_to_gpr[26], preg21_recover_table_to_gpr[26], preg20_recover_table_to_gpr[26],
                                 preg19_recover_table_to_gpr[26], preg18_recover_table_to_gpr[26], preg17_recover_table_to_gpr[26], preg16_recover_table_to_gpr[26],
                                 preg15_recover_table_to_gpr[26], preg14_recover_table_to_gpr[26], preg13_recover_table_to_gpr[26], preg12_recover_table_to_gpr[26],
                                 preg11_recover_table_to_gpr[26], preg10_recover_table_to_gpr[26], preg9_recover_table_to_gpr[26],  preg8_recover_table_to_gpr[26] ,
                                 preg7_recover_table_to_gpr[26],  preg6_recover_table_to_gpr[26],  preg5_recover_table_to_gpr[26],  preg4_recover_table_to_gpr[26] ,
                                 preg3_recover_table_to_gpr[26],  preg2_recover_table_to_gpr[26],  preg1_recover_table_to_gpr[26],  preg0_recover_table_to_gpr[26]};
    assign gpr27_recover_table = {preg63_recover_table_to_gpr[27], preg62_recover_table_to_gpr[27], preg61_recover_table_to_gpr[27], preg60_recover_table_to_gpr[27],
                                 preg59_recover_table_to_gpr[27], preg58_recover_table_to_gpr[27], preg57_recover_table_to_gpr[27], preg56_recover_table_to_gpr[27],
                                 preg55_recover_table_to_gpr[27], preg54_recover_table_to_gpr[27], preg53_recover_table_to_gpr[27], preg52_recover_table_to_gpr[27],
                                 preg51_recover_table_to_gpr[27], preg50_recover_table_to_gpr[27], preg49_recover_table_to_gpr[27], preg48_recover_table_to_gpr[27],
                                 preg47_recover_table_to_gpr[27], preg46_recover_table_to_gpr[27], preg45_recover_table_to_gpr[27], preg44_recover_table_to_gpr[27],
                                 preg43_recover_table_to_gpr[27], preg42_recover_table_to_gpr[27], preg41_recover_table_to_gpr[27], preg40_recover_table_to_gpr[27],
                                 preg39_recover_table_to_gpr[27], preg38_recover_table_to_gpr[27], preg37_recover_table_to_gpr[27], preg36_recover_table_to_gpr[27],
                                 preg35_recover_table_to_gpr[27], preg34_recover_table_to_gpr[27], preg33_recover_table_to_gpr[27], preg32_recover_table_to_gpr[27],
                                 preg31_recover_table_to_gpr[27], preg30_recover_table_to_gpr[27], preg29_recover_table_to_gpr[27], preg28_recover_table_to_gpr[27],
                                 preg27_recover_table_to_gpr[27], preg26_recover_table_to_gpr[27], preg25_recover_table_to_gpr[27], preg24_recover_table_to_gpr[27],
                                 preg23_recover_table_to_gpr[27], preg22_recover_table_to_gpr[27], preg21_recover_table_to_gpr[27], preg20_recover_table_to_gpr[27],
                                 preg19_recover_table_to_gpr[27], preg18_recover_table_to_gpr[27], preg17_recover_table_to_gpr[27], preg16_recover_table_to_gpr[27],
                                 preg15_recover_table_to_gpr[27], preg14_recover_table_to_gpr[27], preg13_recover_table_to_gpr[27], preg12_recover_table_to_gpr[27],
                                 preg11_recover_table_to_gpr[27], preg10_recover_table_to_gpr[27], preg9_recover_table_to_gpr[27],  preg8_recover_table_to_gpr[27] ,
                                 preg7_recover_table_to_gpr[27],  preg6_recover_table_to_gpr[27],  preg5_recover_table_to_gpr[27],  preg4_recover_table_to_gpr[27] ,
                                 preg3_recover_table_to_gpr[27],  preg2_recover_table_to_gpr[27],  preg1_recover_table_to_gpr[27],  preg0_recover_table_to_gpr[27]};
    assign gpr28_recover_table = {preg63_recover_table_to_gpr[28], preg62_recover_table_to_gpr[28], preg61_recover_table_to_gpr[28], preg60_recover_table_to_gpr[28],
                                 preg59_recover_table_to_gpr[28], preg58_recover_table_to_gpr[28], preg57_recover_table_to_gpr[28], preg56_recover_table_to_gpr[28],
                                 preg55_recover_table_to_gpr[28], preg54_recover_table_to_gpr[28], preg53_recover_table_to_gpr[28], preg52_recover_table_to_gpr[28],
                                 preg51_recover_table_to_gpr[28], preg50_recover_table_to_gpr[28], preg49_recover_table_to_gpr[28], preg48_recover_table_to_gpr[28],
                                 preg47_recover_table_to_gpr[28], preg46_recover_table_to_gpr[28], preg45_recover_table_to_gpr[28], preg44_recover_table_to_gpr[28],
                                 preg43_recover_table_to_gpr[28], preg42_recover_table_to_gpr[28], preg41_recover_table_to_gpr[28], preg40_recover_table_to_gpr[28],
                                 preg39_recover_table_to_gpr[28], preg38_recover_table_to_gpr[28], preg37_recover_table_to_gpr[28], preg36_recover_table_to_gpr[28],
                                 preg35_recover_table_to_gpr[28], preg34_recover_table_to_gpr[28], preg33_recover_table_to_gpr[28], preg32_recover_table_to_gpr[28],
                                 preg31_recover_table_to_gpr[28], preg30_recover_table_to_gpr[28], preg29_recover_table_to_gpr[28], preg28_recover_table_to_gpr[28],
                                 preg27_recover_table_to_gpr[28], preg26_recover_table_to_gpr[28], preg25_recover_table_to_gpr[28], preg24_recover_table_to_gpr[28],
                                 preg23_recover_table_to_gpr[28], preg22_recover_table_to_gpr[28], preg21_recover_table_to_gpr[28], preg20_recover_table_to_gpr[28],
                                 preg19_recover_table_to_gpr[28], preg18_recover_table_to_gpr[28], preg17_recover_table_to_gpr[28], preg16_recover_table_to_gpr[28],
                                 preg15_recover_table_to_gpr[28], preg14_recover_table_to_gpr[28], preg13_recover_table_to_gpr[28], preg12_recover_table_to_gpr[28],
                                 preg11_recover_table_to_gpr[28], preg10_recover_table_to_gpr[28], preg9_recover_table_to_gpr[28],  preg8_recover_table_to_gpr[28] ,
                                 preg7_recover_table_to_gpr[28],  preg6_recover_table_to_gpr[28],  preg5_recover_table_to_gpr[28],  preg4_recover_table_to_gpr[28] ,
                                 preg3_recover_table_to_gpr[28],  preg2_recover_table_to_gpr[28],  preg1_recover_table_to_gpr[28],  preg0_recover_table_to_gpr[28]};
    assign gpr29_recover_table = {preg63_recover_table_to_gpr[29], preg62_recover_table_to_gpr[29], preg61_recover_table_to_gpr[29], preg60_recover_table_to_gpr[29],
                                 preg59_recover_table_to_gpr[29], preg58_recover_table_to_gpr[29], preg57_recover_table_to_gpr[29], preg56_recover_table_to_gpr[29],
                                 preg55_recover_table_to_gpr[29], preg54_recover_table_to_gpr[29], preg53_recover_table_to_gpr[29], preg52_recover_table_to_gpr[29],
                                 preg51_recover_table_to_gpr[29], preg50_recover_table_to_gpr[29], preg49_recover_table_to_gpr[29], preg48_recover_table_to_gpr[29],
                                 preg47_recover_table_to_gpr[29], preg46_recover_table_to_gpr[29], preg45_recover_table_to_gpr[29], preg44_recover_table_to_gpr[29],
                                 preg43_recover_table_to_gpr[29], preg42_recover_table_to_gpr[29], preg41_recover_table_to_gpr[29], preg40_recover_table_to_gpr[29],
                                 preg39_recover_table_to_gpr[29], preg38_recover_table_to_gpr[29], preg37_recover_table_to_gpr[29], preg36_recover_table_to_gpr[29],
                                 preg35_recover_table_to_gpr[29], preg34_recover_table_to_gpr[29], preg33_recover_table_to_gpr[29], preg32_recover_table_to_gpr[29],
                                 preg31_recover_table_to_gpr[29], preg30_recover_table_to_gpr[29], preg29_recover_table_to_gpr[29], preg28_recover_table_to_gpr[29],
                                 preg27_recover_table_to_gpr[29], preg26_recover_table_to_gpr[29], preg25_recover_table_to_gpr[29], preg24_recover_table_to_gpr[29],
                                 preg23_recover_table_to_gpr[29], preg22_recover_table_to_gpr[29], preg21_recover_table_to_gpr[29], preg20_recover_table_to_gpr[29],
                                 preg19_recover_table_to_gpr[29], preg18_recover_table_to_gpr[29], preg17_recover_table_to_gpr[29], preg16_recover_table_to_gpr[29],
                                 preg15_recover_table_to_gpr[29], preg14_recover_table_to_gpr[29], preg13_recover_table_to_gpr[29], preg12_recover_table_to_gpr[29],
                                 preg11_recover_table_to_gpr[29], preg10_recover_table_to_gpr[29], preg9_recover_table_to_gpr[29],  preg8_recover_table_to_gpr[29] ,
                                 preg7_recover_table_to_gpr[29],  preg6_recover_table_to_gpr[29],  preg5_recover_table_to_gpr[29],  preg4_recover_table_to_gpr[29] ,
                                 preg3_recover_table_to_gpr[29],  preg2_recover_table_to_gpr[29],  preg1_recover_table_to_gpr[29],  preg0_recover_table_to_gpr[29]};
    assign gpr30_recover_table = {preg63_recover_table_to_gpr[30], preg62_recover_table_to_gpr[30], preg61_recover_table_to_gpr[30], preg60_recover_table_to_gpr[30],
                                 preg59_recover_table_to_gpr[30], preg58_recover_table_to_gpr[30], preg57_recover_table_to_gpr[30], preg56_recover_table_to_gpr[30],
                                 preg55_recover_table_to_gpr[30], preg54_recover_table_to_gpr[30], preg53_recover_table_to_gpr[30], preg52_recover_table_to_gpr[30],
                                 preg51_recover_table_to_gpr[30], preg50_recover_table_to_gpr[30], preg49_recover_table_to_gpr[30], preg48_recover_table_to_gpr[30],
                                 preg47_recover_table_to_gpr[30], preg46_recover_table_to_gpr[30], preg45_recover_table_to_gpr[30], preg44_recover_table_to_gpr[30],
                                 preg43_recover_table_to_gpr[30], preg42_recover_table_to_gpr[30], preg41_recover_table_to_gpr[30], preg40_recover_table_to_gpr[30],
                                 preg39_recover_table_to_gpr[30], preg38_recover_table_to_gpr[30], preg37_recover_table_to_gpr[30], preg36_recover_table_to_gpr[30],
                                 preg35_recover_table_to_gpr[30], preg34_recover_table_to_gpr[30], preg33_recover_table_to_gpr[30], preg32_recover_table_to_gpr[30],
                                 preg31_recover_table_to_gpr[30], preg30_recover_table_to_gpr[30], preg29_recover_table_to_gpr[30], preg28_recover_table_to_gpr[30],
                                 preg27_recover_table_to_gpr[30], preg26_recover_table_to_gpr[30], preg25_recover_table_to_gpr[30], preg24_recover_table_to_gpr[30],
                                 preg23_recover_table_to_gpr[30], preg22_recover_table_to_gpr[30], preg21_recover_table_to_gpr[30], preg20_recover_table_to_gpr[30],
                                 preg19_recover_table_to_gpr[30], preg18_recover_table_to_gpr[30], preg17_recover_table_to_gpr[30], preg16_recover_table_to_gpr[30],
                                 preg15_recover_table_to_gpr[30], preg14_recover_table_to_gpr[30], preg13_recover_table_to_gpr[30], preg12_recover_table_to_gpr[30],
                                 preg11_recover_table_to_gpr[30], preg10_recover_table_to_gpr[30], preg9_recover_table_to_gpr[30],  preg8_recover_table_to_gpr[30] ,
                                 preg7_recover_table_to_gpr[30],  preg6_recover_table_to_gpr[30],  preg5_recover_table_to_gpr[30],  preg4_recover_table_to_gpr[30] ,
                                 preg3_recover_table_to_gpr[30],  preg2_recover_table_to_gpr[30],  preg1_recover_table_to_gpr[30],  preg0_recover_table_to_gpr[30]};
    assign gpr31_recover_table = {preg63_recover_table_to_gpr[31], preg62_recover_table_to_gpr[31], preg61_recover_table_to_gpr[31], preg60_recover_table_to_gpr[31],
                                 preg59_recover_table_to_gpr[31], preg58_recover_table_to_gpr[31], preg57_recover_table_to_gpr[31], preg56_recover_table_to_gpr[31],
                                 preg55_recover_table_to_gpr[31], preg54_recover_table_to_gpr[31], preg53_recover_table_to_gpr[31], preg52_recover_table_to_gpr[31],
                                 preg51_recover_table_to_gpr[31], preg50_recover_table_to_gpr[31], preg49_recover_table_to_gpr[31], preg48_recover_table_to_gpr[31],
                                 preg47_recover_table_to_gpr[31], preg46_recover_table_to_gpr[31], preg45_recover_table_to_gpr[31], preg44_recover_table_to_gpr[31],
                                 preg43_recover_table_to_gpr[31], preg42_recover_table_to_gpr[31], preg41_recover_table_to_gpr[31], preg40_recover_table_to_gpr[31],
                                 preg39_recover_table_to_gpr[31], preg38_recover_table_to_gpr[31], preg37_recover_table_to_gpr[31], preg36_recover_table_to_gpr[31],
                                 preg35_recover_table_to_gpr[31], preg34_recover_table_to_gpr[31], preg33_recover_table_to_gpr[31], preg32_recover_table_to_gpr[31],
                                 preg31_recover_table_to_gpr[31], preg30_recover_table_to_gpr[31], preg29_recover_table_to_gpr[31], preg28_recover_table_to_gpr[31],
                                 preg27_recover_table_to_gpr[31], preg26_recover_table_to_gpr[31], preg25_recover_table_to_gpr[31], preg24_recover_table_to_gpr[31],
                                 preg23_recover_table_to_gpr[31], preg22_recover_table_to_gpr[31], preg21_recover_table_to_gpr[31], preg20_recover_table_to_gpr[31],
                                 preg19_recover_table_to_gpr[31], preg18_recover_table_to_gpr[31], preg17_recover_table_to_gpr[31], preg16_recover_table_to_gpr[31],
                                 preg15_recover_table_to_gpr[31], preg14_recover_table_to_gpr[31], preg13_recover_table_to_gpr[31], preg12_recover_table_to_gpr[31],
                                 preg11_recover_table_to_gpr[31], preg10_recover_table_to_gpr[31], preg9_recover_table_to_gpr[31],  preg8_recover_table_to_gpr[31] ,
                                 preg7_recover_table_to_gpr[31],  preg6_recover_table_to_gpr[31],  preg5_recover_table_to_gpr[31],  preg4_recover_table_to_gpr[31] ,
                                 preg3_recover_table_to_gpr[31],  preg2_recover_table_to_gpr[31],  preg1_recover_table_to_gpr[31],  preg0_recover_table_to_gpr[31]};
    assign gpr0_recover_mapped  = {6{gpr0_recover_table[0]}}  & 6'd0
                                | {6{gpr0_recover_table[1]}}  & 6'd1
                                | {6{gpr0_recover_table[2]}}  & 6'd2
                                | {6{gpr0_recover_table[3]}}  & 6'd3
                                | {6{gpr0_recover_table[4]}}  & 6'd4
                                | {6{gpr0_recover_table[5]}}  & 6'd5
                                | {6{gpr0_recover_table[6]}}  & 6'd6
                                | {6{gpr0_recover_table[7]}}  & 6'd7
                                | {6{gpr0_recover_table[8]}}  & 6'd8
                                | {6{gpr0_recover_table[9]}}  & 6'd9
                                | {6{gpr0_recover_table[10]}} & 6'd10
                                | {6{gpr0_recover_table[11]}} & 6'd11
                                | {6{gpr0_recover_table[12]}} & 6'd12
                                | {6{gpr0_recover_table[13]}} & 6'd13
                                | {6{gpr0_recover_table[14]}} & 6'd14
                                | {6{gpr0_recover_table[15]}} & 6'd15
                                | {6{gpr0_recover_table[16]}} & 6'd16
                                | {6{gpr0_recover_table[17]}} & 6'd17
                                | {6{gpr0_recover_table[18]}} & 6'd18
                                | {6{gpr0_recover_table[19]}} & 6'd19
                                | {6{gpr0_recover_table[20]}} & 6'd20
                                | {6{gpr0_recover_table[21]}} & 6'd21
                                | {6{gpr0_recover_table[22]}} & 6'd22
                                | {6{gpr0_recover_table[23]}} & 6'd23
                                | {6{gpr0_recover_table[24]}} & 6'd24
                                | {6{gpr0_recover_table[25]}} & 6'd25
                                | {6{gpr0_recover_table[26]}} & 6'd26
                                | {6{gpr0_recover_table[27]}} & 6'd27
                                | {6{gpr0_recover_table[28]}} & 6'd28
                                | {6{gpr0_recover_table[29]}} & 6'd29
                                | {6{gpr0_recover_table[30]}} & 6'd30
                                | {6{gpr0_recover_table[31]}} & 6'd31
                                | {6{gpr0_recover_table[32]}} & 6'd32
                                | {6{gpr0_recover_table[33]}} & 6'd33
                                | {6{gpr0_recover_table[34]}} & 6'd34
                                | {6{gpr0_recover_table[35]}} & 6'd35
                                | {6{gpr0_recover_table[36]}} & 6'd36
                                | {6{gpr0_recover_table[37]}} & 6'd37
                                | {6{gpr0_recover_table[38]}} & 6'd38
                                | {6{gpr0_recover_table[39]}} & 6'd39
                                | {6{gpr0_recover_table[40]}} & 6'd40
                                | {6{gpr0_recover_table[41]}} & 6'd41
                                | {6{gpr0_recover_table[42]}} & 6'd42
                                | {6{gpr0_recover_table[43]}} & 6'd43
                                | {6{gpr0_recover_table[44]}} & 6'd44
                                | {6{gpr0_recover_table[45]}} & 6'd45
                                | {6{gpr0_recover_table[46]}} & 6'd46
                                | {6{gpr0_recover_table[47]}} & 6'd47
                                | {6{gpr0_recover_table[48]}} & 6'd48
                                | {6{gpr0_recover_table[49]}} & 6'd49
                                | {6{gpr0_recover_table[50]}} & 6'd50
                                | {6{gpr0_recover_table[51]}} & 6'd51
                                | {6{gpr0_recover_table[52]}} & 6'd52
                                | {6{gpr0_recover_table[53]}} & 6'd53
                                | {6{gpr0_recover_table[54]}} & 6'd54
                                | {6{gpr0_recover_table[55]}} & 6'd55
                                | {6{gpr0_recover_table[56]}} & 6'd56
                                | {6{gpr0_recover_table[57]}} & 6'd57
                                | {6{gpr0_recover_table[58]}} & 6'd58
                                | {6{gpr0_recover_table[59]}} & 6'd59
                                | {6{gpr0_recover_table[60]}} & 6'd60
                                | {6{gpr0_recover_table[61]}} & 6'd61
                                | {6{gpr0_recover_table[62]}} & 6'd62
                                | {6{gpr0_recover_table[63]}} & 6'd63;
    assign gpr1_recover_mapped  = {6{gpr1_recover_table[0]}}  & 6'd0
                                | {6{gpr1_recover_table[1]}}  & 6'd1
                                | {6{gpr1_recover_table[2]}}  & 6'd2
                                | {6{gpr1_recover_table[3]}}  & 6'd3
                                | {6{gpr1_recover_table[4]}}  & 6'd4
                                | {6{gpr1_recover_table[5]}}  & 6'd5
                                | {6{gpr1_recover_table[6]}}  & 6'd6
                                | {6{gpr1_recover_table[7]}}  & 6'd7
                                | {6{gpr1_recover_table[8]}}  & 6'd8
                                | {6{gpr1_recover_table[9]}}  & 6'd9
                                | {6{gpr1_recover_table[10]}} & 6'd10
                                | {6{gpr1_recover_table[11]}} & 6'd11
                                | {6{gpr1_recover_table[12]}} & 6'd12
                                | {6{gpr1_recover_table[13]}} & 6'd13
                                | {6{gpr1_recover_table[14]}} & 6'd14
                                | {6{gpr1_recover_table[15]}} & 6'd15
                                | {6{gpr1_recover_table[16]}} & 6'd16
                                | {6{gpr1_recover_table[17]}} & 6'd17
                                | {6{gpr1_recover_table[18]}} & 6'd18
                                | {6{gpr1_recover_table[19]}} & 6'd19
                                | {6{gpr1_recover_table[20]}} & 6'd20
                                | {6{gpr1_recover_table[21]}} & 6'd21
                                | {6{gpr1_recover_table[22]}} & 6'd22
                                | {6{gpr1_recover_table[23]}} & 6'd23
                                | {6{gpr1_recover_table[24]}} & 6'd24
                                | {6{gpr1_recover_table[25]}} & 6'd25
                                | {6{gpr1_recover_table[26]}} & 6'd26
                                | {6{gpr1_recover_table[27]}} & 6'd27
                                | {6{gpr1_recover_table[28]}} & 6'd28
                                | {6{gpr1_recover_table[29]}} & 6'd29
                                | {6{gpr1_recover_table[30]}} & 6'd30
                                | {6{gpr1_recover_table[31]}} & 6'd31
                                | {6{gpr1_recover_table[32]}} & 6'd32
                                | {6{gpr1_recover_table[33]}} & 6'd33
                                | {6{gpr1_recover_table[34]}} & 6'd34
                                | {6{gpr1_recover_table[35]}} & 6'd35
                                | {6{gpr1_recover_table[36]}} & 6'd36
                                | {6{gpr1_recover_table[37]}} & 6'd37
                                | {6{gpr1_recover_table[38]}} & 6'd38
                                | {6{gpr1_recover_table[39]}} & 6'd39
                                | {6{gpr1_recover_table[40]}} & 6'd40
                                | {6{gpr1_recover_table[41]}} & 6'd41
                                | {6{gpr1_recover_table[42]}} & 6'd42
                                | {6{gpr1_recover_table[43]}} & 6'd43
                                | {6{gpr1_recover_table[44]}} & 6'd44
                                | {6{gpr1_recover_table[45]}} & 6'd45
                                | {6{gpr1_recover_table[46]}} & 6'd46
                                | {6{gpr1_recover_table[47]}} & 6'd47
                                | {6{gpr1_recover_table[48]}} & 6'd48
                                | {6{gpr1_recover_table[49]}} & 6'd49
                                | {6{gpr1_recover_table[50]}} & 6'd50
                                | {6{gpr1_recover_table[51]}} & 6'd51
                                | {6{gpr1_recover_table[52]}} & 6'd52
                                | {6{gpr1_recover_table[53]}} & 6'd53
                                | {6{gpr1_recover_table[54]}} & 6'd54
                                | {6{gpr1_recover_table[55]}} & 6'd55
                                | {6{gpr1_recover_table[56]}} & 6'd56
                                | {6{gpr1_recover_table[57]}} & 6'd57
                                | {6{gpr1_recover_table[58]}} & 6'd58
                                | {6{gpr1_recover_table[59]}} & 6'd59
                                | {6{gpr1_recover_table[60]}} & 6'd60
                                | {6{gpr1_recover_table[61]}} & 6'd61
                                | {6{gpr1_recover_table[62]}} & 6'd62
                                | {6{gpr1_recover_table[63]}} & 6'd63;
    assign gpr2_recover_mapped  = {6{gpr2_recover_table[0]}}  & 6'd0
                                | {6{gpr2_recover_table[1]}}  & 6'd1
                                | {6{gpr2_recover_table[2]}}  & 6'd2
                                | {6{gpr2_recover_table[3]}}  & 6'd3
                                | {6{gpr2_recover_table[4]}}  & 6'd4
                                | {6{gpr2_recover_table[5]}}  & 6'd5
                                | {6{gpr2_recover_table[6]}}  & 6'd6
                                | {6{gpr2_recover_table[7]}}  & 6'd7
                                | {6{gpr2_recover_table[8]}}  & 6'd8
                                | {6{gpr2_recover_table[9]}}  & 6'd9
                                | {6{gpr2_recover_table[10]}} & 6'd10
                                | {6{gpr2_recover_table[11]}} & 6'd11
                                | {6{gpr2_recover_table[12]}} & 6'd12
                                | {6{gpr2_recover_table[13]}} & 6'd13
                                | {6{gpr2_recover_table[14]}} & 6'd14
                                | {6{gpr2_recover_table[15]}} & 6'd15
                                | {6{gpr2_recover_table[16]}} & 6'd16
                                | {6{gpr2_recover_table[17]}} & 6'd17
                                | {6{gpr2_recover_table[18]}} & 6'd18
                                | {6{gpr2_recover_table[19]}} & 6'd19
                                | {6{gpr2_recover_table[20]}} & 6'd20
                                | {6{gpr2_recover_table[21]}} & 6'd21
                                | {6{gpr2_recover_table[22]}} & 6'd22
                                | {6{gpr2_recover_table[23]}} & 6'd23
                                | {6{gpr2_recover_table[24]}} & 6'd24
                                | {6{gpr2_recover_table[25]}} & 6'd25
                                | {6{gpr2_recover_table[26]}} & 6'd26
                                | {6{gpr2_recover_table[27]}} & 6'd27
                                | {6{gpr2_recover_table[28]}} & 6'd28
                                | {6{gpr2_recover_table[29]}} & 6'd29
                                | {6{gpr2_recover_table[30]}} & 6'd30
                                | {6{gpr2_recover_table[31]}} & 6'd31
                                | {6{gpr2_recover_table[32]}} & 6'd32
                                | {6{gpr2_recover_table[33]}} & 6'd33
                                | {6{gpr2_recover_table[34]}} & 6'd34
                                | {6{gpr2_recover_table[35]}} & 6'd35
                                | {6{gpr2_recover_table[36]}} & 6'd36
                                | {6{gpr2_recover_table[37]}} & 6'd37
                                | {6{gpr2_recover_table[38]}} & 6'd38
                                | {6{gpr2_recover_table[39]}} & 6'd39
                                | {6{gpr2_recover_table[40]}} & 6'd40
                                | {6{gpr2_recover_table[41]}} & 6'd41
                                | {6{gpr2_recover_table[42]}} & 6'd42
                                | {6{gpr2_recover_table[43]}} & 6'd43
                                | {6{gpr2_recover_table[44]}} & 6'd44
                                | {6{gpr2_recover_table[45]}} & 6'd45
                                | {6{gpr2_recover_table[46]}} & 6'd46
                                | {6{gpr2_recover_table[47]}} & 6'd47
                                | {6{gpr2_recover_table[48]}} & 6'd48
                                | {6{gpr2_recover_table[49]}} & 6'd49
                                | {6{gpr2_recover_table[50]}} & 6'd50
                                | {6{gpr2_recover_table[51]}} & 6'd51
                                | {6{gpr2_recover_table[52]}} & 6'd52
                                | {6{gpr2_recover_table[53]}} & 6'd53
                                | {6{gpr2_recover_table[54]}} & 6'd54
                                | {6{gpr2_recover_table[55]}} & 6'd55
                                | {6{gpr2_recover_table[56]}} & 6'd56
                                | {6{gpr2_recover_table[57]}} & 6'd57
                                | {6{gpr2_recover_table[58]}} & 6'd58
                                | {6{gpr2_recover_table[59]}} & 6'd59
                                | {6{gpr2_recover_table[60]}} & 6'd60
                                | {6{gpr2_recover_table[61]}} & 6'd61
                                | {6{gpr2_recover_table[62]}} & 6'd62
                                | {6{gpr2_recover_table[63]}} & 6'd63;
    assign gpr3_recover_mapped  = {6{gpr3_recover_table[0]}}  & 6'd0
                                | {6{gpr3_recover_table[1]}}  & 6'd1
                                | {6{gpr3_recover_table[2]}}  & 6'd2
                                | {6{gpr3_recover_table[3]}}  & 6'd3
                                | {6{gpr3_recover_table[4]}}  & 6'd4
                                | {6{gpr3_recover_table[5]}}  & 6'd5
                                | {6{gpr3_recover_table[6]}}  & 6'd6
                                | {6{gpr3_recover_table[7]}}  & 6'd7
                                | {6{gpr3_recover_table[8]}}  & 6'd8
                                | {6{gpr3_recover_table[9]}}  & 6'd9
                                | {6{gpr3_recover_table[10]}} & 6'd10
                                | {6{gpr3_recover_table[11]}} & 6'd11
                                | {6{gpr3_recover_table[12]}} & 6'd12
                                | {6{gpr3_recover_table[13]}} & 6'd13
                                | {6{gpr3_recover_table[14]}} & 6'd14
                                | {6{gpr3_recover_table[15]}} & 6'd15
                                | {6{gpr3_recover_table[16]}} & 6'd16
                                | {6{gpr3_recover_table[17]}} & 6'd17
                                | {6{gpr3_recover_table[18]}} & 6'd18
                                | {6{gpr3_recover_table[19]}} & 6'd19
                                | {6{gpr3_recover_table[20]}} & 6'd20
                                | {6{gpr3_recover_table[21]}} & 6'd21
                                | {6{gpr3_recover_table[22]}} & 6'd22
                                | {6{gpr3_recover_table[23]}} & 6'd23
                                | {6{gpr3_recover_table[24]}} & 6'd24
                                | {6{gpr3_recover_table[25]}} & 6'd25
                                | {6{gpr3_recover_table[26]}} & 6'd26
                                | {6{gpr3_recover_table[27]}} & 6'd27
                                | {6{gpr3_recover_table[28]}} & 6'd28
                                | {6{gpr3_recover_table[29]}} & 6'd29
                                | {6{gpr3_recover_table[30]}} & 6'd30
                                | {6{gpr3_recover_table[31]}} & 6'd31
                                | {6{gpr3_recover_table[32]}} & 6'd32
                                | {6{gpr3_recover_table[33]}} & 6'd33
                                | {6{gpr3_recover_table[34]}} & 6'd34
                                | {6{gpr3_recover_table[35]}} & 6'd35
                                | {6{gpr3_recover_table[36]}} & 6'd36
                                | {6{gpr3_recover_table[37]}} & 6'd37
                                | {6{gpr3_recover_table[38]}} & 6'd38
                                | {6{gpr3_recover_table[39]}} & 6'd39
                                | {6{gpr3_recover_table[40]}} & 6'd40
                                | {6{gpr3_recover_table[41]}} & 6'd41
                                | {6{gpr3_recover_table[42]}} & 6'd42
                                | {6{gpr3_recover_table[43]}} & 6'd43
                                | {6{gpr3_recover_table[44]}} & 6'd44
                                | {6{gpr3_recover_table[45]}} & 6'd45
                                | {6{gpr3_recover_table[46]}} & 6'd46
                                | {6{gpr3_recover_table[47]}} & 6'd47
                                | {6{gpr3_recover_table[48]}} & 6'd48
                                | {6{gpr3_recover_table[49]}} & 6'd49
                                | {6{gpr3_recover_table[50]}} & 6'd50
                                | {6{gpr3_recover_table[51]}} & 6'd51
                                | {6{gpr3_recover_table[52]}} & 6'd52
                                | {6{gpr3_recover_table[53]}} & 6'd53
                                | {6{gpr3_recover_table[54]}} & 6'd54
                                | {6{gpr3_recover_table[55]}} & 6'd55
                                | {6{gpr3_recover_table[56]}} & 6'd56
                                | {6{gpr3_recover_table[57]}} & 6'd57
                                | {6{gpr3_recover_table[58]}} & 6'd58
                                | {6{gpr3_recover_table[59]}} & 6'd59
                                | {6{gpr3_recover_table[60]}} & 6'd60
                                | {6{gpr3_recover_table[61]}} & 6'd61
                                | {6{gpr3_recover_table[62]}} & 6'd62
                                | {6{gpr3_recover_table[63]}} & 6'd63;
    assign gpr4_recover_mapped  = {6{gpr4_recover_table[0]}}  & 6'd0
                                | {6{gpr4_recover_table[1]}}  & 6'd1
                                | {6{gpr4_recover_table[2]}}  & 6'd2
                                | {6{gpr4_recover_table[3]}}  & 6'd3
                                | {6{gpr4_recover_table[4]}}  & 6'd4
                                | {6{gpr4_recover_table[5]}}  & 6'd5
                                | {6{gpr4_recover_table[6]}}  & 6'd6
                                | {6{gpr4_recover_table[7]}}  & 6'd7
                                | {6{gpr4_recover_table[8]}}  & 6'd8
                                | {6{gpr4_recover_table[9]}}  & 6'd9
                                | {6{gpr4_recover_table[10]}} & 6'd10
                                | {6{gpr4_recover_table[11]}} & 6'd11
                                | {6{gpr4_recover_table[12]}} & 6'd12
                                | {6{gpr4_recover_table[13]}} & 6'd13
                                | {6{gpr4_recover_table[14]}} & 6'd14
                                | {6{gpr4_recover_table[15]}} & 6'd15
                                | {6{gpr4_recover_table[16]}} & 6'd16
                                | {6{gpr4_recover_table[17]}} & 6'd17
                                | {6{gpr4_recover_table[18]}} & 6'd18
                                | {6{gpr4_recover_table[19]}} & 6'd19
                                | {6{gpr4_recover_table[20]}} & 6'd20
                                | {6{gpr4_recover_table[21]}} & 6'd21
                                | {6{gpr4_recover_table[22]}} & 6'd22
                                | {6{gpr4_recover_table[23]}} & 6'd23
                                | {6{gpr4_recover_table[24]}} & 6'd24
                                | {6{gpr4_recover_table[25]}} & 6'd25
                                | {6{gpr4_recover_table[26]}} & 6'd26
                                | {6{gpr4_recover_table[27]}} & 6'd27
                                | {6{gpr4_recover_table[28]}} & 6'd28
                                | {6{gpr4_recover_table[29]}} & 6'd29
                                | {6{gpr4_recover_table[30]}} & 6'd30
                                | {6{gpr4_recover_table[31]}} & 6'd31
                                | {6{gpr4_recover_table[32]}} & 6'd32
                                | {6{gpr4_recover_table[33]}} & 6'd33
                                | {6{gpr4_recover_table[34]}} & 6'd34
                                | {6{gpr4_recover_table[35]}} & 6'd35
                                | {6{gpr4_recover_table[36]}} & 6'd36
                                | {6{gpr4_recover_table[37]}} & 6'd37
                                | {6{gpr4_recover_table[38]}} & 6'd38
                                | {6{gpr4_recover_table[39]}} & 6'd39
                                | {6{gpr4_recover_table[40]}} & 6'd40
                                | {6{gpr4_recover_table[41]}} & 6'd41
                                | {6{gpr4_recover_table[42]}} & 6'd42
                                | {6{gpr4_recover_table[43]}} & 6'd43
                                | {6{gpr4_recover_table[44]}} & 6'd44
                                | {6{gpr4_recover_table[45]}} & 6'd45
                                | {6{gpr4_recover_table[46]}} & 6'd46
                                | {6{gpr4_recover_table[47]}} & 6'd47
                                | {6{gpr4_recover_table[48]}} & 6'd48
                                | {6{gpr4_recover_table[49]}} & 6'd49
                                | {6{gpr4_recover_table[50]}} & 6'd50
                                | {6{gpr4_recover_table[51]}} & 6'd51
                                | {6{gpr4_recover_table[52]}} & 6'd52
                                | {6{gpr4_recover_table[53]}} & 6'd53
                                | {6{gpr4_recover_table[54]}} & 6'd54
                                | {6{gpr4_recover_table[55]}} & 6'd55
                                | {6{gpr4_recover_table[56]}} & 6'd56
                                | {6{gpr4_recover_table[57]}} & 6'd57
                                | {6{gpr4_recover_table[58]}} & 6'd58
                                | {6{gpr4_recover_table[59]}} & 6'd59
                                | {6{gpr4_recover_table[60]}} & 6'd60
                                | {6{gpr4_recover_table[61]}} & 6'd61
                                | {6{gpr4_recover_table[62]}} & 6'd62
                                | {6{gpr4_recover_table[63]}} & 6'd63;
    assign gpr5_recover_mapped  = {6{gpr5_recover_table[0]}}  & 6'd0
                                | {6{gpr5_recover_table[1]}}  & 6'd1
                                | {6{gpr5_recover_table[2]}}  & 6'd2
                                | {6{gpr5_recover_table[3]}}  & 6'd3
                                | {6{gpr5_recover_table[4]}}  & 6'd4
                                | {6{gpr5_recover_table[5]}}  & 6'd5
                                | {6{gpr5_recover_table[6]}}  & 6'd6
                                | {6{gpr5_recover_table[7]}}  & 6'd7
                                | {6{gpr5_recover_table[8]}}  & 6'd8
                                | {6{gpr5_recover_table[9]}}  & 6'd9
                                | {6{gpr5_recover_table[10]}} & 6'd10
                                | {6{gpr5_recover_table[11]}} & 6'd11
                                | {6{gpr5_recover_table[12]}} & 6'd12
                                | {6{gpr5_recover_table[13]}} & 6'd13
                                | {6{gpr5_recover_table[14]}} & 6'd14
                                | {6{gpr5_recover_table[15]}} & 6'd15
                                | {6{gpr5_recover_table[16]}} & 6'd16
                                | {6{gpr5_recover_table[17]}} & 6'd17
                                | {6{gpr5_recover_table[18]}} & 6'd18
                                | {6{gpr5_recover_table[19]}} & 6'd19
                                | {6{gpr5_recover_table[20]}} & 6'd20
                                | {6{gpr5_recover_table[21]}} & 6'd21
                                | {6{gpr5_recover_table[22]}} & 6'd22
                                | {6{gpr5_recover_table[23]}} & 6'd23
                                | {6{gpr5_recover_table[24]}} & 6'd24
                                | {6{gpr5_recover_table[25]}} & 6'd25
                                | {6{gpr5_recover_table[26]}} & 6'd26
                                | {6{gpr5_recover_table[27]}} & 6'd27
                                | {6{gpr5_recover_table[28]}} & 6'd28
                                | {6{gpr5_recover_table[29]}} & 6'd29
                                | {6{gpr5_recover_table[30]}} & 6'd30
                                | {6{gpr5_recover_table[31]}} & 6'd31
                                | {6{gpr5_recover_table[32]}} & 6'd32
                                | {6{gpr5_recover_table[33]}} & 6'd33
                                | {6{gpr5_recover_table[34]}} & 6'd34
                                | {6{gpr5_recover_table[35]}} & 6'd35
                                | {6{gpr5_recover_table[36]}} & 6'd36
                                | {6{gpr5_recover_table[37]}} & 6'd37
                                | {6{gpr5_recover_table[38]}} & 6'd38
                                | {6{gpr5_recover_table[39]}} & 6'd39
                                | {6{gpr5_recover_table[40]}} & 6'd40
                                | {6{gpr5_recover_table[41]}} & 6'd41
                                | {6{gpr5_recover_table[42]}} & 6'd42
                                | {6{gpr5_recover_table[43]}} & 6'd43
                                | {6{gpr5_recover_table[44]}} & 6'd44
                                | {6{gpr5_recover_table[45]}} & 6'd45
                                | {6{gpr5_recover_table[46]}} & 6'd46
                                | {6{gpr5_recover_table[47]}} & 6'd47
                                | {6{gpr5_recover_table[48]}} & 6'd48
                                | {6{gpr5_recover_table[49]}} & 6'd49
                                | {6{gpr5_recover_table[50]}} & 6'd50
                                | {6{gpr5_recover_table[51]}} & 6'd51
                                | {6{gpr5_recover_table[52]}} & 6'd52
                                | {6{gpr5_recover_table[53]}} & 6'd53
                                | {6{gpr5_recover_table[54]}} & 6'd54
                                | {6{gpr5_recover_table[55]}} & 6'd55
                                | {6{gpr5_recover_table[56]}} & 6'd56
                                | {6{gpr5_recover_table[57]}} & 6'd57
                                | {6{gpr5_recover_table[58]}} & 6'd58
                                | {6{gpr5_recover_table[59]}} & 6'd59
                                | {6{gpr5_recover_table[60]}} & 6'd60
                                | {6{gpr5_recover_table[61]}} & 6'd61
                                | {6{gpr5_recover_table[62]}} & 6'd62
                                | {6{gpr5_recover_table[63]}} & 6'd63;
    assign gpr6_recover_mapped  = {6{gpr6_recover_table[0]}}  & 6'd0
                                | {6{gpr6_recover_table[1]}}  & 6'd1
                                | {6{gpr6_recover_table[2]}}  & 6'd2
                                | {6{gpr6_recover_table[3]}}  & 6'd3
                                | {6{gpr6_recover_table[4]}}  & 6'd4
                                | {6{gpr6_recover_table[5]}}  & 6'd5
                                | {6{gpr6_recover_table[6]}}  & 6'd6
                                | {6{gpr6_recover_table[7]}}  & 6'd7
                                | {6{gpr6_recover_table[8]}}  & 6'd8
                                | {6{gpr6_recover_table[9]}}  & 6'd9
                                | {6{gpr6_recover_table[10]}} & 6'd10
                                | {6{gpr6_recover_table[11]}} & 6'd11
                                | {6{gpr6_recover_table[12]}} & 6'd12
                                | {6{gpr6_recover_table[13]}} & 6'd13
                                | {6{gpr6_recover_table[14]}} & 6'd14
                                | {6{gpr6_recover_table[15]}} & 6'd15
                                | {6{gpr6_recover_table[16]}} & 6'd16
                                | {6{gpr6_recover_table[17]}} & 6'd17
                                | {6{gpr6_recover_table[18]}} & 6'd18
                                | {6{gpr6_recover_table[19]}} & 6'd19
                                | {6{gpr6_recover_table[20]}} & 6'd20
                                | {6{gpr6_recover_table[21]}} & 6'd21
                                | {6{gpr6_recover_table[22]}} & 6'd22
                                | {6{gpr6_recover_table[23]}} & 6'd23
                                | {6{gpr6_recover_table[24]}} & 6'd24
                                | {6{gpr6_recover_table[25]}} & 6'd25
                                | {6{gpr6_recover_table[26]}} & 6'd26
                                | {6{gpr6_recover_table[27]}} & 6'd27
                                | {6{gpr6_recover_table[28]}} & 6'd28
                                | {6{gpr6_recover_table[29]}} & 6'd29
                                | {6{gpr6_recover_table[30]}} & 6'd30
                                | {6{gpr6_recover_table[31]}} & 6'd31
                                | {6{gpr6_recover_table[32]}} & 6'd32
                                | {6{gpr6_recover_table[33]}} & 6'd33
                                | {6{gpr6_recover_table[34]}} & 6'd34
                                | {6{gpr6_recover_table[35]}} & 6'd35
                                | {6{gpr6_recover_table[36]}} & 6'd36
                                | {6{gpr6_recover_table[37]}} & 6'd37
                                | {6{gpr6_recover_table[38]}} & 6'd38
                                | {6{gpr6_recover_table[39]}} & 6'd39
                                | {6{gpr6_recover_table[40]}} & 6'd40
                                | {6{gpr6_recover_table[41]}} & 6'd41
                                | {6{gpr6_recover_table[42]}} & 6'd42
                                | {6{gpr6_recover_table[43]}} & 6'd43
                                | {6{gpr6_recover_table[44]}} & 6'd44
                                | {6{gpr6_recover_table[45]}} & 6'd45
                                | {6{gpr6_recover_table[46]}} & 6'd46
                                | {6{gpr6_recover_table[47]}} & 6'd47
                                | {6{gpr6_recover_table[48]}} & 6'd48
                                | {6{gpr6_recover_table[49]}} & 6'd49
                                | {6{gpr6_recover_table[50]}} & 6'd50
                                | {6{gpr6_recover_table[51]}} & 6'd51
                                | {6{gpr6_recover_table[52]}} & 6'd52
                                | {6{gpr6_recover_table[53]}} & 6'd53
                                | {6{gpr6_recover_table[54]}} & 6'd54
                                | {6{gpr6_recover_table[55]}} & 6'd55
                                | {6{gpr6_recover_table[56]}} & 6'd56
                                | {6{gpr6_recover_table[57]}} & 6'd57
                                | {6{gpr6_recover_table[58]}} & 6'd58
                                | {6{gpr6_recover_table[59]}} & 6'd59
                                | {6{gpr6_recover_table[60]}} & 6'd60
                                | {6{gpr6_recover_table[61]}} & 6'd61
                                | {6{gpr6_recover_table[62]}} & 6'd62
                                | {6{gpr6_recover_table[63]}} & 6'd63;
    assign gpr7_recover_mapped  = {6{gpr7_recover_table[0]}}  & 6'd0
                                | {6{gpr7_recover_table[1]}}  & 6'd1
                                | {6{gpr7_recover_table[2]}}  & 6'd2
                                | {6{gpr7_recover_table[3]}}  & 6'd3
                                | {6{gpr7_recover_table[4]}}  & 6'd4
                                | {6{gpr7_recover_table[5]}}  & 6'd5
                                | {6{gpr7_recover_table[6]}}  & 6'd6
                                | {6{gpr7_recover_table[7]}}  & 6'd7
                                | {6{gpr7_recover_table[8]}}  & 6'd8
                                | {6{gpr7_recover_table[9]}}  & 6'd9
                                | {6{gpr7_recover_table[10]}} & 6'd10
                                | {6{gpr7_recover_table[11]}} & 6'd11
                                | {6{gpr7_recover_table[12]}} & 6'd12
                                | {6{gpr7_recover_table[13]}} & 6'd13
                                | {6{gpr7_recover_table[14]}} & 6'd14
                                | {6{gpr7_recover_table[15]}} & 6'd15
                                | {6{gpr7_recover_table[16]}} & 6'd16
                                | {6{gpr7_recover_table[17]}} & 6'd17
                                | {6{gpr7_recover_table[18]}} & 6'd18
                                | {6{gpr7_recover_table[19]}} & 6'd19
                                | {6{gpr7_recover_table[20]}} & 6'd20
                                | {6{gpr7_recover_table[21]}} & 6'd21
                                | {6{gpr7_recover_table[22]}} & 6'd22
                                | {6{gpr7_recover_table[23]}} & 6'd23
                                | {6{gpr7_recover_table[24]}} & 6'd24
                                | {6{gpr7_recover_table[25]}} & 6'd25
                                | {6{gpr7_recover_table[26]}} & 6'd26
                                | {6{gpr7_recover_table[27]}} & 6'd27
                                | {6{gpr7_recover_table[28]}} & 6'd28
                                | {6{gpr7_recover_table[29]}} & 6'd29
                                | {6{gpr7_recover_table[30]}} & 6'd30
                                | {6{gpr7_recover_table[31]}} & 6'd31
                                | {6{gpr7_recover_table[32]}} & 6'd32
                                | {6{gpr7_recover_table[33]}} & 6'd33
                                | {6{gpr7_recover_table[34]}} & 6'd34
                                | {6{gpr7_recover_table[35]}} & 6'd35
                                | {6{gpr7_recover_table[36]}} & 6'd36
                                | {6{gpr7_recover_table[37]}} & 6'd37
                                | {6{gpr7_recover_table[38]}} & 6'd38
                                | {6{gpr7_recover_table[39]}} & 6'd39
                                | {6{gpr7_recover_table[40]}} & 6'd40
                                | {6{gpr7_recover_table[41]}} & 6'd41
                                | {6{gpr7_recover_table[42]}} & 6'd42
                                | {6{gpr7_recover_table[43]}} & 6'd43
                                | {6{gpr7_recover_table[44]}} & 6'd44
                                | {6{gpr7_recover_table[45]}} & 6'd45
                                | {6{gpr7_recover_table[46]}} & 6'd46
                                | {6{gpr7_recover_table[47]}} & 6'd47
                                | {6{gpr7_recover_table[48]}} & 6'd48
                                | {6{gpr7_recover_table[49]}} & 6'd49
                                | {6{gpr7_recover_table[50]}} & 6'd50
                                | {6{gpr7_recover_table[51]}} & 6'd51
                                | {6{gpr7_recover_table[52]}} & 6'd52
                                | {6{gpr7_recover_table[53]}} & 6'd53
                                | {6{gpr7_recover_table[54]}} & 6'd54
                                | {6{gpr7_recover_table[55]}} & 6'd55
                                | {6{gpr7_recover_table[56]}} & 6'd56
                                | {6{gpr7_recover_table[57]}} & 6'd57
                                | {6{gpr7_recover_table[58]}} & 6'd58
                                | {6{gpr7_recover_table[59]}} & 6'd59
                                | {6{gpr7_recover_table[60]}} & 6'd60
                                | {6{gpr7_recover_table[61]}} & 6'd61
                                | {6{gpr7_recover_table[62]}} & 6'd62
                                | {6{gpr7_recover_table[63]}} & 6'd63;
    assign gpr8_recover_mapped  = {6{gpr8_recover_table[0]}}  & 6'd0
                                | {6{gpr8_recover_table[1]}}  & 6'd1
                                | {6{gpr8_recover_table[2]}}  & 6'd2
                                | {6{gpr8_recover_table[3]}}  & 6'd3
                                | {6{gpr8_recover_table[4]}}  & 6'd4
                                | {6{gpr8_recover_table[5]}}  & 6'd5
                                | {6{gpr8_recover_table[6]}}  & 6'd6
                                | {6{gpr8_recover_table[7]}}  & 6'd7
                                | {6{gpr8_recover_table[8]}}  & 6'd8
                                | {6{gpr8_recover_table[9]}}  & 6'd9
                                | {6{gpr8_recover_table[10]}} & 6'd10
                                | {6{gpr8_recover_table[11]}} & 6'd11
                                | {6{gpr8_recover_table[12]}} & 6'd12
                                | {6{gpr8_recover_table[13]}} & 6'd13
                                | {6{gpr8_recover_table[14]}} & 6'd14
                                | {6{gpr8_recover_table[15]}} & 6'd15
                                | {6{gpr8_recover_table[16]}} & 6'd16
                                | {6{gpr8_recover_table[17]}} & 6'd17
                                | {6{gpr8_recover_table[18]}} & 6'd18
                                | {6{gpr8_recover_table[19]}} & 6'd19
                                | {6{gpr8_recover_table[20]}} & 6'd20
                                | {6{gpr8_recover_table[21]}} & 6'd21
                                | {6{gpr8_recover_table[22]}} & 6'd22
                                | {6{gpr8_recover_table[23]}} & 6'd23
                                | {6{gpr8_recover_table[24]}} & 6'd24
                                | {6{gpr8_recover_table[25]}} & 6'd25
                                | {6{gpr8_recover_table[26]}} & 6'd26
                                | {6{gpr8_recover_table[27]}} & 6'd27
                                | {6{gpr8_recover_table[28]}} & 6'd28
                                | {6{gpr8_recover_table[29]}} & 6'd29
                                | {6{gpr8_recover_table[30]}} & 6'd30
                                | {6{gpr8_recover_table[31]}} & 6'd31
                                | {6{gpr8_recover_table[32]}} & 6'd32
                                | {6{gpr8_recover_table[33]}} & 6'd33
                                | {6{gpr8_recover_table[34]}} & 6'd34
                                | {6{gpr8_recover_table[35]}} & 6'd35
                                | {6{gpr8_recover_table[36]}} & 6'd36
                                | {6{gpr8_recover_table[37]}} & 6'd37
                                | {6{gpr8_recover_table[38]}} & 6'd38
                                | {6{gpr8_recover_table[39]}} & 6'd39
                                | {6{gpr8_recover_table[40]}} & 6'd40
                                | {6{gpr8_recover_table[41]}} & 6'd41
                                | {6{gpr8_recover_table[42]}} & 6'd42
                                | {6{gpr8_recover_table[43]}} & 6'd43
                                | {6{gpr8_recover_table[44]}} & 6'd44
                                | {6{gpr8_recover_table[45]}} & 6'd45
                                | {6{gpr8_recover_table[46]}} & 6'd46
                                | {6{gpr8_recover_table[47]}} & 6'd47
                                | {6{gpr8_recover_table[48]}} & 6'd48
                                | {6{gpr8_recover_table[49]}} & 6'd49
                                | {6{gpr8_recover_table[50]}} & 6'd50
                                | {6{gpr8_recover_table[51]}} & 6'd51
                                | {6{gpr8_recover_table[52]}} & 6'd52
                                | {6{gpr8_recover_table[53]}} & 6'd53
                                | {6{gpr8_recover_table[54]}} & 6'd54
                                | {6{gpr8_recover_table[55]}} & 6'd55
                                | {6{gpr8_recover_table[56]}} & 6'd56
                                | {6{gpr8_recover_table[57]}} & 6'd57
                                | {6{gpr8_recover_table[58]}} & 6'd58
                                | {6{gpr8_recover_table[59]}} & 6'd59
                                | {6{gpr8_recover_table[60]}} & 6'd60
                                | {6{gpr8_recover_table[61]}} & 6'd61
                                | {6{gpr8_recover_table[62]}} & 6'd62
                                | {6{gpr8_recover_table[63]}} & 6'd63;
    assign gpr9_recover_mapped  = {6{gpr9_recover_table[0]}}  & 6'd0
                                | {6{gpr9_recover_table[1]}}  & 6'd1
                                | {6{gpr9_recover_table[2]}}  & 6'd2
                                | {6{gpr9_recover_table[3]}}  & 6'd3
                                | {6{gpr9_recover_table[4]}}  & 6'd4
                                | {6{gpr9_recover_table[5]}}  & 6'd5
                                | {6{gpr9_recover_table[6]}}  & 6'd6
                                | {6{gpr9_recover_table[7]}}  & 6'd7
                                | {6{gpr9_recover_table[8]}}  & 6'd8
                                | {6{gpr9_recover_table[9]}}  & 6'd9
                                | {6{gpr9_recover_table[10]}} & 6'd10
                                | {6{gpr9_recover_table[11]}} & 6'd11
                                | {6{gpr9_recover_table[12]}} & 6'd12
                                | {6{gpr9_recover_table[13]}} & 6'd13
                                | {6{gpr9_recover_table[14]}} & 6'd14
                                | {6{gpr9_recover_table[15]}} & 6'd15
                                | {6{gpr9_recover_table[16]}} & 6'd16
                                | {6{gpr9_recover_table[17]}} & 6'd17
                                | {6{gpr9_recover_table[18]}} & 6'd18
                                | {6{gpr9_recover_table[19]}} & 6'd19
                                | {6{gpr9_recover_table[20]}} & 6'd20
                                | {6{gpr9_recover_table[21]}} & 6'd21
                                | {6{gpr9_recover_table[22]}} & 6'd22
                                | {6{gpr9_recover_table[23]}} & 6'd23
                                | {6{gpr9_recover_table[24]}} & 6'd24
                                | {6{gpr9_recover_table[25]}} & 6'd25
                                | {6{gpr9_recover_table[26]}} & 6'd26
                                | {6{gpr9_recover_table[27]}} & 6'd27
                                | {6{gpr9_recover_table[28]}} & 6'd28
                                | {6{gpr9_recover_table[29]}} & 6'd29
                                | {6{gpr9_recover_table[30]}} & 6'd30
                                | {6{gpr9_recover_table[31]}} & 6'd31
                                | {6{gpr9_recover_table[32]}} & 6'd32
                                | {6{gpr9_recover_table[33]}} & 6'd33
                                | {6{gpr9_recover_table[34]}} & 6'd34
                                | {6{gpr9_recover_table[35]}} & 6'd35
                                | {6{gpr9_recover_table[36]}} & 6'd36
                                | {6{gpr9_recover_table[37]}} & 6'd37
                                | {6{gpr9_recover_table[38]}} & 6'd38
                                | {6{gpr9_recover_table[39]}} & 6'd39
                                | {6{gpr9_recover_table[40]}} & 6'd40
                                | {6{gpr9_recover_table[41]}} & 6'd41
                                | {6{gpr9_recover_table[42]}} & 6'd42
                                | {6{gpr9_recover_table[43]}} & 6'd43
                                | {6{gpr9_recover_table[44]}} & 6'd44
                                | {6{gpr9_recover_table[45]}} & 6'd45
                                | {6{gpr9_recover_table[46]}} & 6'd46
                                | {6{gpr9_recover_table[47]}} & 6'd47
                                | {6{gpr9_recover_table[48]}} & 6'd48
                                | {6{gpr9_recover_table[49]}} & 6'd49
                                | {6{gpr9_recover_table[50]}} & 6'd50
                                | {6{gpr9_recover_table[51]}} & 6'd51
                                | {6{gpr9_recover_table[52]}} & 6'd52
                                | {6{gpr9_recover_table[53]}} & 6'd53
                                | {6{gpr9_recover_table[54]}} & 6'd54
                                | {6{gpr9_recover_table[55]}} & 6'd55
                                | {6{gpr9_recover_table[56]}} & 6'd56
                                | {6{gpr9_recover_table[57]}} & 6'd57
                                | {6{gpr9_recover_table[58]}} & 6'd58
                                | {6{gpr9_recover_table[59]}} & 6'd59
                                | {6{gpr9_recover_table[60]}} & 6'd60
                                | {6{gpr9_recover_table[61]}} & 6'd61
                                | {6{gpr9_recover_table[62]}} & 6'd62
                                | {6{gpr9_recover_table[63]}} & 6'd63;
    assign gpr10_recover_mapped = {6{gpr10_recover_table[0]}}  & 6'd0
                                | {6{gpr10_recover_table[1]}}  & 6'd1
                                | {6{gpr10_recover_table[2]}}  & 6'd2
                                | {6{gpr10_recover_table[3]}}  & 6'd3
                                | {6{gpr10_recover_table[4]}}  & 6'd4
                                | {6{gpr10_recover_table[5]}}  & 6'd5
                                | {6{gpr10_recover_table[6]}}  & 6'd6
                                | {6{gpr10_recover_table[7]}}  & 6'd7
                                | {6{gpr10_recover_table[8]}}  & 6'd8
                                | {6{gpr10_recover_table[9]}}  & 6'd9
                                | {6{gpr10_recover_table[10]}} & 6'd10
                                | {6{gpr10_recover_table[11]}} & 6'd11
                                | {6{gpr10_recover_table[12]}} & 6'd12
                                | {6{gpr10_recover_table[13]}} & 6'd13
                                | {6{gpr10_recover_table[14]}} & 6'd14
                                | {6{gpr10_recover_table[15]}} & 6'd15
                                | {6{gpr10_recover_table[16]}} & 6'd16
                                | {6{gpr10_recover_table[17]}} & 6'd17
                                | {6{gpr10_recover_table[18]}} & 6'd18
                                | {6{gpr10_recover_table[19]}} & 6'd19
                                | {6{gpr10_recover_table[20]}} & 6'd20
                                | {6{gpr10_recover_table[21]}} & 6'd21
                                | {6{gpr10_recover_table[22]}} & 6'd22
                                | {6{gpr10_recover_table[23]}} & 6'd23
                                | {6{gpr10_recover_table[24]}} & 6'd24
                                | {6{gpr10_recover_table[25]}} & 6'd25
                                | {6{gpr10_recover_table[26]}} & 6'd26
                                | {6{gpr10_recover_table[27]}} & 6'd27
                                | {6{gpr10_recover_table[28]}} & 6'd28
                                | {6{gpr10_recover_table[29]}} & 6'd29
                                | {6{gpr10_recover_table[30]}} & 6'd30
                                | {6{gpr10_recover_table[31]}} & 6'd31
                                | {6{gpr10_recover_table[32]}} & 6'd32
                                | {6{gpr10_recover_table[33]}} & 6'd33
                                | {6{gpr10_recover_table[34]}} & 6'd34
                                | {6{gpr10_recover_table[35]}} & 6'd35
                                | {6{gpr10_recover_table[36]}} & 6'd36
                                | {6{gpr10_recover_table[37]}} & 6'd37
                                | {6{gpr10_recover_table[38]}} & 6'd38
                                | {6{gpr10_recover_table[39]}} & 6'd39
                                | {6{gpr10_recover_table[40]}} & 6'd40
                                | {6{gpr10_recover_table[41]}} & 6'd41
                                | {6{gpr10_recover_table[42]}} & 6'd42
                                | {6{gpr10_recover_table[43]}} & 6'd43
                                | {6{gpr10_recover_table[44]}} & 6'd44
                                | {6{gpr10_recover_table[45]}} & 6'd45
                                | {6{gpr10_recover_table[46]}} & 6'd46
                                | {6{gpr10_recover_table[47]}} & 6'd47
                                | {6{gpr10_recover_table[48]}} & 6'd48
                                | {6{gpr10_recover_table[49]}} & 6'd49
                                | {6{gpr10_recover_table[50]}} & 6'd50
                                | {6{gpr10_recover_table[51]}} & 6'd51
                                | {6{gpr10_recover_table[52]}} & 6'd52
                                | {6{gpr10_recover_table[53]}} & 6'd53
                                | {6{gpr10_recover_table[54]}} & 6'd54
                                | {6{gpr10_recover_table[55]}} & 6'd55
                                | {6{gpr10_recover_table[56]}} & 6'd56
                                | {6{gpr10_recover_table[57]}} & 6'd57
                                | {6{gpr10_recover_table[58]}} & 6'd58
                                | {6{gpr10_recover_table[59]}} & 6'd59
                                | {6{gpr10_recover_table[60]}} & 6'd60
                                | {6{gpr10_recover_table[61]}} & 6'd61
                                | {6{gpr10_recover_table[62]}} & 6'd62
                                | {6{gpr10_recover_table[63]}} & 6'd63;
    assign gpr11_recover_mapped = {6{gpr11_recover_table[0]}}  & 6'd0
                                | {6{gpr11_recover_table[1]}}  & 6'd1
                                | {6{gpr11_recover_table[2]}}  & 6'd2
                                | {6{gpr11_recover_table[3]}}  & 6'd3
                                | {6{gpr11_recover_table[4]}}  & 6'd4
                                | {6{gpr11_recover_table[5]}}  & 6'd5
                                | {6{gpr11_recover_table[6]}}  & 6'd6
                                | {6{gpr11_recover_table[7]}}  & 6'd7
                                | {6{gpr11_recover_table[8]}}  & 6'd8
                                | {6{gpr11_recover_table[9]}}  & 6'd9
                                | {6{gpr11_recover_table[10]}} & 6'd10
                                | {6{gpr11_recover_table[11]}} & 6'd11
                                | {6{gpr11_recover_table[12]}} & 6'd12
                                | {6{gpr11_recover_table[13]}} & 6'd13
                                | {6{gpr11_recover_table[14]}} & 6'd14
                                | {6{gpr11_recover_table[15]}} & 6'd15
                                | {6{gpr11_recover_table[16]}} & 6'd16
                                | {6{gpr11_recover_table[17]}} & 6'd17
                                | {6{gpr11_recover_table[18]}} & 6'd18
                                | {6{gpr11_recover_table[19]}} & 6'd19
                                | {6{gpr11_recover_table[20]}} & 6'd20
                                | {6{gpr11_recover_table[21]}} & 6'd21
                                | {6{gpr11_recover_table[22]}} & 6'd22
                                | {6{gpr11_recover_table[23]}} & 6'd23
                                | {6{gpr11_recover_table[24]}} & 6'd24
                                | {6{gpr11_recover_table[25]}} & 6'd25
                                | {6{gpr11_recover_table[26]}} & 6'd26
                                | {6{gpr11_recover_table[27]}} & 6'd27
                                | {6{gpr11_recover_table[28]}} & 6'd28
                                | {6{gpr11_recover_table[29]}} & 6'd29
                                | {6{gpr11_recover_table[30]}} & 6'd30
                                | {6{gpr11_recover_table[31]}} & 6'd31
                                | {6{gpr11_recover_table[32]}} & 6'd32
                                | {6{gpr11_recover_table[33]}} & 6'd33
                                | {6{gpr11_recover_table[34]}} & 6'd34
                                | {6{gpr11_recover_table[35]}} & 6'd35
                                | {6{gpr11_recover_table[36]}} & 6'd36
                                | {6{gpr11_recover_table[37]}} & 6'd37
                                | {6{gpr11_recover_table[38]}} & 6'd38
                                | {6{gpr11_recover_table[39]}} & 6'd39
                                | {6{gpr11_recover_table[40]}} & 6'd40
                                | {6{gpr11_recover_table[41]}} & 6'd41
                                | {6{gpr11_recover_table[42]}} & 6'd42
                                | {6{gpr11_recover_table[43]}} & 6'd43
                                | {6{gpr11_recover_table[44]}} & 6'd44
                                | {6{gpr11_recover_table[45]}} & 6'd45
                                | {6{gpr11_recover_table[46]}} & 6'd46
                                | {6{gpr11_recover_table[47]}} & 6'd47
                                | {6{gpr11_recover_table[48]}} & 6'd48
                                | {6{gpr11_recover_table[49]}} & 6'd49
                                | {6{gpr11_recover_table[50]}} & 6'd50
                                | {6{gpr11_recover_table[51]}} & 6'd51
                                | {6{gpr11_recover_table[52]}} & 6'd52
                                | {6{gpr11_recover_table[53]}} & 6'd53
                                | {6{gpr11_recover_table[54]}} & 6'd54
                                | {6{gpr11_recover_table[55]}} & 6'd55
                                | {6{gpr11_recover_table[56]}} & 6'd56
                                | {6{gpr11_recover_table[57]}} & 6'd57
                                | {6{gpr11_recover_table[58]}} & 6'd58
                                | {6{gpr11_recover_table[59]}} & 6'd59
                                | {6{gpr11_recover_table[60]}} & 6'd60
                                | {6{gpr11_recover_table[61]}} & 6'd61
                                | {6{gpr11_recover_table[62]}} & 6'd62
                                | {6{gpr11_recover_table[63]}} & 6'd63;
    assign gpr12_recover_mapped = {6{gpr12_recover_table[0]}}  & 6'd0
                                | {6{gpr12_recover_table[1]}}  & 6'd1
                                | {6{gpr12_recover_table[2]}}  & 6'd2
                                | {6{gpr12_recover_table[3]}}  & 6'd3
                                | {6{gpr12_recover_table[4]}}  & 6'd4
                                | {6{gpr12_recover_table[5]}}  & 6'd5
                                | {6{gpr12_recover_table[6]}}  & 6'd6
                                | {6{gpr12_recover_table[7]}}  & 6'd7
                                | {6{gpr12_recover_table[8]}}  & 6'd8
                                | {6{gpr12_recover_table[9]}}  & 6'd9
                                | {6{gpr12_recover_table[10]}} & 6'd10
                                | {6{gpr12_recover_table[11]}} & 6'd11
                                | {6{gpr12_recover_table[12]}} & 6'd12
                                | {6{gpr12_recover_table[13]}} & 6'd13
                                | {6{gpr12_recover_table[14]}} & 6'd14
                                | {6{gpr12_recover_table[15]}} & 6'd15
                                | {6{gpr12_recover_table[16]}} & 6'd16
                                | {6{gpr12_recover_table[17]}} & 6'd17
                                | {6{gpr12_recover_table[18]}} & 6'd18
                                | {6{gpr12_recover_table[19]}} & 6'd19
                                | {6{gpr12_recover_table[20]}} & 6'd20
                                | {6{gpr12_recover_table[21]}} & 6'd21
                                | {6{gpr12_recover_table[22]}} & 6'd22
                                | {6{gpr12_recover_table[23]}} & 6'd23
                                | {6{gpr12_recover_table[24]}} & 6'd24
                                | {6{gpr12_recover_table[25]}} & 6'd25
                                | {6{gpr12_recover_table[26]}} & 6'd26
                                | {6{gpr12_recover_table[27]}} & 6'd27
                                | {6{gpr12_recover_table[28]}} & 6'd28
                                | {6{gpr12_recover_table[29]}} & 6'd29
                                | {6{gpr12_recover_table[30]}} & 6'd30
                                | {6{gpr12_recover_table[31]}} & 6'd31
                                | {6{gpr12_recover_table[32]}} & 6'd32
                                | {6{gpr12_recover_table[33]}} & 6'd33
                                | {6{gpr12_recover_table[34]}} & 6'd34
                                | {6{gpr12_recover_table[35]}} & 6'd35
                                | {6{gpr12_recover_table[36]}} & 6'd36
                                | {6{gpr12_recover_table[37]}} & 6'd37
                                | {6{gpr12_recover_table[38]}} & 6'd38
                                | {6{gpr12_recover_table[39]}} & 6'd39
                                | {6{gpr12_recover_table[40]}} & 6'd40
                                | {6{gpr12_recover_table[41]}} & 6'd41
                                | {6{gpr12_recover_table[42]}} & 6'd42
                                | {6{gpr12_recover_table[43]}} & 6'd43
                                | {6{gpr12_recover_table[44]}} & 6'd44
                                | {6{gpr12_recover_table[45]}} & 6'd45
                                | {6{gpr12_recover_table[46]}} & 6'd46
                                | {6{gpr12_recover_table[47]}} & 6'd47
                                | {6{gpr12_recover_table[48]}} & 6'd48
                                | {6{gpr12_recover_table[49]}} & 6'd49
                                | {6{gpr12_recover_table[50]}} & 6'd50
                                | {6{gpr12_recover_table[51]}} & 6'd51
                                | {6{gpr12_recover_table[52]}} & 6'd52
                                | {6{gpr12_recover_table[53]}} & 6'd53
                                | {6{gpr12_recover_table[54]}} & 6'd54
                                | {6{gpr12_recover_table[55]}} & 6'd55
                                | {6{gpr12_recover_table[56]}} & 6'd56
                                | {6{gpr12_recover_table[57]}} & 6'd57
                                | {6{gpr12_recover_table[58]}} & 6'd58
                                | {6{gpr12_recover_table[59]}} & 6'd59
                                | {6{gpr12_recover_table[60]}} & 6'd60
                                | {6{gpr12_recover_table[61]}} & 6'd61
                                | {6{gpr12_recover_table[62]}} & 6'd62
                                | {6{gpr12_recover_table[63]}} & 6'd63;
    assign gpr13_recover_mapped = {6{gpr13_recover_table[0]}}  & 6'd0
                                | {6{gpr13_recover_table[1]}}  & 6'd1
                                | {6{gpr13_recover_table[2]}}  & 6'd2
                                | {6{gpr13_recover_table[3]}}  & 6'd3
                                | {6{gpr13_recover_table[4]}}  & 6'd4
                                | {6{gpr13_recover_table[5]}}  & 6'd5
                                | {6{gpr13_recover_table[6]}}  & 6'd6
                                | {6{gpr13_recover_table[7]}}  & 6'd7
                                | {6{gpr13_recover_table[8]}}  & 6'd8
                                | {6{gpr13_recover_table[9]}}  & 6'd9
                                | {6{gpr13_recover_table[10]}} & 6'd10
                                | {6{gpr13_recover_table[11]}} & 6'd11
                                | {6{gpr13_recover_table[12]}} & 6'd12
                                | {6{gpr13_recover_table[13]}} & 6'd13
                                | {6{gpr13_recover_table[14]}} & 6'd14
                                | {6{gpr13_recover_table[15]}} & 6'd15
                                | {6{gpr13_recover_table[16]}} & 6'd16
                                | {6{gpr13_recover_table[17]}} & 6'd17
                                | {6{gpr13_recover_table[18]}} & 6'd18
                                | {6{gpr13_recover_table[19]}} & 6'd19
                                | {6{gpr13_recover_table[20]}} & 6'd20
                                | {6{gpr13_recover_table[21]}} & 6'd21
                                | {6{gpr13_recover_table[22]}} & 6'd22
                                | {6{gpr13_recover_table[23]}} & 6'd23
                                | {6{gpr13_recover_table[24]}} & 6'd24
                                | {6{gpr13_recover_table[25]}} & 6'd25
                                | {6{gpr13_recover_table[26]}} & 6'd26
                                | {6{gpr13_recover_table[27]}} & 6'd27
                                | {6{gpr13_recover_table[28]}} & 6'd28
                                | {6{gpr13_recover_table[29]}} & 6'd29
                                | {6{gpr13_recover_table[30]}} & 6'd30
                                | {6{gpr13_recover_table[31]}} & 6'd31
                                | {6{gpr13_recover_table[32]}} & 6'd32
                                | {6{gpr13_recover_table[33]}} & 6'd33
                                | {6{gpr13_recover_table[34]}} & 6'd34
                                | {6{gpr13_recover_table[35]}} & 6'd35
                                | {6{gpr13_recover_table[36]}} & 6'd36
                                | {6{gpr13_recover_table[37]}} & 6'd37
                                | {6{gpr13_recover_table[38]}} & 6'd38
                                | {6{gpr13_recover_table[39]}} & 6'd39
                                | {6{gpr13_recover_table[40]}} & 6'd40
                                | {6{gpr13_recover_table[41]}} & 6'd41
                                | {6{gpr13_recover_table[42]}} & 6'd42
                                | {6{gpr13_recover_table[43]}} & 6'd43
                                | {6{gpr13_recover_table[44]}} & 6'd44
                                | {6{gpr13_recover_table[45]}} & 6'd45
                                | {6{gpr13_recover_table[46]}} & 6'd46
                                | {6{gpr13_recover_table[47]}} & 6'd47
                                | {6{gpr13_recover_table[48]}} & 6'd48
                                | {6{gpr13_recover_table[49]}} & 6'd49
                                | {6{gpr13_recover_table[50]}} & 6'd50
                                | {6{gpr13_recover_table[51]}} & 6'd51
                                | {6{gpr13_recover_table[52]}} & 6'd52
                                | {6{gpr13_recover_table[53]}} & 6'd53
                                | {6{gpr13_recover_table[54]}} & 6'd54
                                | {6{gpr13_recover_table[55]}} & 6'd55
                                | {6{gpr13_recover_table[56]}} & 6'd56
                                | {6{gpr13_recover_table[57]}} & 6'd57
                                | {6{gpr13_recover_table[58]}} & 6'd58
                                | {6{gpr13_recover_table[59]}} & 6'd59
                                | {6{gpr13_recover_table[60]}} & 6'd60
                                | {6{gpr13_recover_table[61]}} & 6'd61
                                | {6{gpr13_recover_table[62]}} & 6'd62
                                | {6{gpr13_recover_table[63]}} & 6'd63;
    assign gpr14_recover_mapped = {6{gpr14_recover_table[0]}}  & 6'd0
                                | {6{gpr14_recover_table[1]}}  & 6'd1
                                | {6{gpr14_recover_table[2]}}  & 6'd2
                                | {6{gpr14_recover_table[3]}}  & 6'd3
                                | {6{gpr14_recover_table[4]}}  & 6'd4
                                | {6{gpr14_recover_table[5]}}  & 6'd5
                                | {6{gpr14_recover_table[6]}}  & 6'd6
                                | {6{gpr14_recover_table[7]}}  & 6'd7
                                | {6{gpr14_recover_table[8]}}  & 6'd8
                                | {6{gpr14_recover_table[9]}}  & 6'd9
                                | {6{gpr14_recover_table[10]}} & 6'd10
                                | {6{gpr14_recover_table[11]}} & 6'd11
                                | {6{gpr14_recover_table[12]}} & 6'd12
                                | {6{gpr14_recover_table[13]}} & 6'd13
                                | {6{gpr14_recover_table[14]}} & 6'd14
                                | {6{gpr14_recover_table[15]}} & 6'd15
                                | {6{gpr14_recover_table[16]}} & 6'd16
                                | {6{gpr14_recover_table[17]}} & 6'd17
                                | {6{gpr14_recover_table[18]}} & 6'd18
                                | {6{gpr14_recover_table[19]}} & 6'd19
                                | {6{gpr14_recover_table[20]}} & 6'd20
                                | {6{gpr14_recover_table[21]}} & 6'd21
                                | {6{gpr14_recover_table[22]}} & 6'd22
                                | {6{gpr14_recover_table[23]}} & 6'd23
                                | {6{gpr14_recover_table[24]}} & 6'd24
                                | {6{gpr14_recover_table[25]}} & 6'd25
                                | {6{gpr14_recover_table[26]}} & 6'd26
                                | {6{gpr14_recover_table[27]}} & 6'd27
                                | {6{gpr14_recover_table[28]}} & 6'd28
                                | {6{gpr14_recover_table[29]}} & 6'd29
                                | {6{gpr14_recover_table[30]}} & 6'd30
                                | {6{gpr14_recover_table[31]}} & 6'd31
                                | {6{gpr14_recover_table[32]}} & 6'd32
                                | {6{gpr14_recover_table[33]}} & 6'd33
                                | {6{gpr14_recover_table[34]}} & 6'd34
                                | {6{gpr14_recover_table[35]}} & 6'd35
                                | {6{gpr14_recover_table[36]}} & 6'd36
                                | {6{gpr14_recover_table[37]}} & 6'd37
                                | {6{gpr14_recover_table[38]}} & 6'd38
                                | {6{gpr14_recover_table[39]}} & 6'd39
                                | {6{gpr14_recover_table[40]}} & 6'd40
                                | {6{gpr14_recover_table[41]}} & 6'd41
                                | {6{gpr14_recover_table[42]}} & 6'd42
                                | {6{gpr14_recover_table[43]}} & 6'd43
                                | {6{gpr14_recover_table[44]}} & 6'd44
                                | {6{gpr14_recover_table[45]}} & 6'd45
                                | {6{gpr14_recover_table[46]}} & 6'd46
                                | {6{gpr14_recover_table[47]}} & 6'd47
                                | {6{gpr14_recover_table[48]}} & 6'd48
                                | {6{gpr14_recover_table[49]}} & 6'd49
                                | {6{gpr14_recover_table[50]}} & 6'd50
                                | {6{gpr14_recover_table[51]}} & 6'd51
                                | {6{gpr14_recover_table[52]}} & 6'd52
                                | {6{gpr14_recover_table[53]}} & 6'd53
                                | {6{gpr14_recover_table[54]}} & 6'd54
                                | {6{gpr14_recover_table[55]}} & 6'd55
                                | {6{gpr14_recover_table[56]}} & 6'd56
                                | {6{gpr14_recover_table[57]}} & 6'd57
                                | {6{gpr14_recover_table[58]}} & 6'd58
                                | {6{gpr14_recover_table[59]}} & 6'd59
                                | {6{gpr14_recover_table[60]}} & 6'd60
                                | {6{gpr14_recover_table[61]}} & 6'd61
                                | {6{gpr14_recover_table[62]}} & 6'd62
                                | {6{gpr14_recover_table[63]}} & 6'd63;
    assign gpr15_recover_mapped = {6{gpr15_recover_table[0]}}  & 6'd0
                                | {6{gpr15_recover_table[1]}}  & 6'd1
                                | {6{gpr15_recover_table[2]}}  & 6'd2
                                | {6{gpr15_recover_table[3]}}  & 6'd3
                                | {6{gpr15_recover_table[4]}}  & 6'd4
                                | {6{gpr15_recover_table[5]}}  & 6'd5
                                | {6{gpr15_recover_table[6]}}  & 6'd6
                                | {6{gpr15_recover_table[7]}}  & 6'd7
                                | {6{gpr15_recover_table[8]}}  & 6'd8
                                | {6{gpr15_recover_table[9]}}  & 6'd9
                                | {6{gpr15_recover_table[10]}} & 6'd10
                                | {6{gpr15_recover_table[11]}} & 6'd11
                                | {6{gpr15_recover_table[12]}} & 6'd12
                                | {6{gpr15_recover_table[13]}} & 6'd13
                                | {6{gpr15_recover_table[14]}} & 6'd14
                                | {6{gpr15_recover_table[15]}} & 6'd15
                                | {6{gpr15_recover_table[16]}} & 6'd16
                                | {6{gpr15_recover_table[17]}} & 6'd17
                                | {6{gpr15_recover_table[18]}} & 6'd18
                                | {6{gpr15_recover_table[19]}} & 6'd19
                                | {6{gpr15_recover_table[20]}} & 6'd20
                                | {6{gpr15_recover_table[21]}} & 6'd21
                                | {6{gpr15_recover_table[22]}} & 6'd22
                                | {6{gpr15_recover_table[23]}} & 6'd23
                                | {6{gpr15_recover_table[24]}} & 6'd24
                                | {6{gpr15_recover_table[25]}} & 6'd25
                                | {6{gpr15_recover_table[26]}} & 6'd26
                                | {6{gpr15_recover_table[27]}} & 6'd27
                                | {6{gpr15_recover_table[28]}} & 6'd28
                                | {6{gpr15_recover_table[29]}} & 6'd29
                                | {6{gpr15_recover_table[30]}} & 6'd30
                                | {6{gpr15_recover_table[31]}} & 6'd31
                                | {6{gpr15_recover_table[32]}} & 6'd32
                                | {6{gpr15_recover_table[33]}} & 6'd33
                                | {6{gpr15_recover_table[34]}} & 6'd34
                                | {6{gpr15_recover_table[35]}} & 6'd35
                                | {6{gpr15_recover_table[36]}} & 6'd36
                                | {6{gpr15_recover_table[37]}} & 6'd37
                                | {6{gpr15_recover_table[38]}} & 6'd38
                                | {6{gpr15_recover_table[39]}} & 6'd39
                                | {6{gpr15_recover_table[40]}} & 6'd40
                                | {6{gpr15_recover_table[41]}} & 6'd41
                                | {6{gpr15_recover_table[42]}} & 6'd42
                                | {6{gpr15_recover_table[43]}} & 6'd43
                                | {6{gpr15_recover_table[44]}} & 6'd44
                                | {6{gpr15_recover_table[45]}} & 6'd45
                                | {6{gpr15_recover_table[46]}} & 6'd46
                                | {6{gpr15_recover_table[47]}} & 6'd47
                                | {6{gpr15_recover_table[48]}} & 6'd48
                                | {6{gpr15_recover_table[49]}} & 6'd49
                                | {6{gpr15_recover_table[50]}} & 6'd50
                                | {6{gpr15_recover_table[51]}} & 6'd51
                                | {6{gpr15_recover_table[52]}} & 6'd52
                                | {6{gpr15_recover_table[53]}} & 6'd53
                                | {6{gpr15_recover_table[54]}} & 6'd54
                                | {6{gpr15_recover_table[55]}} & 6'd55
                                | {6{gpr15_recover_table[56]}} & 6'd56
                                | {6{gpr15_recover_table[57]}} & 6'd57
                                | {6{gpr15_recover_table[58]}} & 6'd58
                                | {6{gpr15_recover_table[59]}} & 6'd59
                                | {6{gpr15_recover_table[60]}} & 6'd60
                                | {6{gpr15_recover_table[61]}} & 6'd61
                                | {6{gpr15_recover_table[62]}} & 6'd62
                                | {6{gpr15_recover_table[63]}} & 6'd63;
    assign gpr16_recover_mapped = {6{gpr16_recover_table[0]}}  & 6'd0
                                | {6{gpr16_recover_table[1]}}  & 6'd1
                                | {6{gpr16_recover_table[2]}}  & 6'd2
                                | {6{gpr16_recover_table[3]}}  & 6'd3
                                | {6{gpr16_recover_table[4]}}  & 6'd4
                                | {6{gpr16_recover_table[5]}}  & 6'd5
                                | {6{gpr16_recover_table[6]}}  & 6'd6
                                | {6{gpr16_recover_table[7]}}  & 6'd7
                                | {6{gpr16_recover_table[8]}}  & 6'd8
                                | {6{gpr16_recover_table[9]}}  & 6'd9
                                | {6{gpr16_recover_table[10]}} & 6'd10
                                | {6{gpr16_recover_table[11]}} & 6'd11
                                | {6{gpr16_recover_table[12]}} & 6'd12
                                | {6{gpr16_recover_table[13]}} & 6'd13
                                | {6{gpr16_recover_table[14]}} & 6'd14
                                | {6{gpr16_recover_table[15]}} & 6'd15
                                | {6{gpr16_recover_table[16]}} & 6'd16
                                | {6{gpr16_recover_table[17]}} & 6'd17
                                | {6{gpr16_recover_table[18]}} & 6'd18
                                | {6{gpr16_recover_table[19]}} & 6'd19
                                | {6{gpr16_recover_table[20]}} & 6'd20
                                | {6{gpr16_recover_table[21]}} & 6'd21
                                | {6{gpr16_recover_table[22]}} & 6'd22
                                | {6{gpr16_recover_table[23]}} & 6'd23
                                | {6{gpr16_recover_table[24]}} & 6'd24
                                | {6{gpr16_recover_table[25]}} & 6'd25
                                | {6{gpr16_recover_table[26]}} & 6'd26
                                | {6{gpr16_recover_table[27]}} & 6'd27
                                | {6{gpr16_recover_table[28]}} & 6'd28
                                | {6{gpr16_recover_table[29]}} & 6'd29
                                | {6{gpr16_recover_table[30]}} & 6'd30
                                | {6{gpr16_recover_table[31]}} & 6'd31
                                | {6{gpr16_recover_table[32]}} & 6'd32
                                | {6{gpr16_recover_table[33]}} & 6'd33
                                | {6{gpr16_recover_table[34]}} & 6'd34
                                | {6{gpr16_recover_table[35]}} & 6'd35
                                | {6{gpr16_recover_table[36]}} & 6'd36
                                | {6{gpr16_recover_table[37]}} & 6'd37
                                | {6{gpr16_recover_table[38]}} & 6'd38
                                | {6{gpr16_recover_table[39]}} & 6'd39
                                | {6{gpr16_recover_table[40]}} & 6'd40
                                | {6{gpr16_recover_table[41]}} & 6'd41
                                | {6{gpr16_recover_table[42]}} & 6'd42
                                | {6{gpr16_recover_table[43]}} & 6'd43
                                | {6{gpr16_recover_table[44]}} & 6'd44
                                | {6{gpr16_recover_table[45]}} & 6'd45
                                | {6{gpr16_recover_table[46]}} & 6'd46
                                | {6{gpr16_recover_table[47]}} & 6'd47
                                | {6{gpr16_recover_table[48]}} & 6'd48
                                | {6{gpr16_recover_table[49]}} & 6'd49
                                | {6{gpr16_recover_table[50]}} & 6'd50
                                | {6{gpr16_recover_table[51]}} & 6'd51
                                | {6{gpr16_recover_table[52]}} & 6'd52
                                | {6{gpr16_recover_table[53]}} & 6'd53
                                | {6{gpr16_recover_table[54]}} & 6'd54
                                | {6{gpr16_recover_table[55]}} & 6'd55
                                | {6{gpr16_recover_table[56]}} & 6'd56
                                | {6{gpr16_recover_table[57]}} & 6'd57
                                | {6{gpr16_recover_table[58]}} & 6'd58
                                | {6{gpr16_recover_table[59]}} & 6'd59
                                | {6{gpr16_recover_table[60]}} & 6'd60
                                | {6{gpr16_recover_table[61]}} & 6'd61
                                | {6{gpr16_recover_table[62]}} & 6'd62
                                | {6{gpr16_recover_table[63]}} & 6'd63;
    assign gpr17_recover_mapped = {6{gpr17_recover_table[0]}}  & 6'd0
                                | {6{gpr17_recover_table[1]}}  & 6'd1
                                | {6{gpr17_recover_table[2]}}  & 6'd2
                                | {6{gpr17_recover_table[3]}}  & 6'd3
                                | {6{gpr17_recover_table[4]}}  & 6'd4
                                | {6{gpr17_recover_table[5]}}  & 6'd5
                                | {6{gpr17_recover_table[6]}}  & 6'd6
                                | {6{gpr17_recover_table[7]}}  & 6'd7
                                | {6{gpr17_recover_table[8]}}  & 6'd8
                                | {6{gpr17_recover_table[9]}}  & 6'd9
                                | {6{gpr17_recover_table[10]}} & 6'd10
                                | {6{gpr17_recover_table[11]}} & 6'd11
                                | {6{gpr17_recover_table[12]}} & 6'd12
                                | {6{gpr17_recover_table[13]}} & 6'd13
                                | {6{gpr17_recover_table[14]}} & 6'd14
                                | {6{gpr17_recover_table[15]}} & 6'd15
                                | {6{gpr17_recover_table[16]}} & 6'd16
                                | {6{gpr17_recover_table[17]}} & 6'd17
                                | {6{gpr17_recover_table[18]}} & 6'd18
                                | {6{gpr17_recover_table[19]}} & 6'd19
                                | {6{gpr17_recover_table[20]}} & 6'd20
                                | {6{gpr17_recover_table[21]}} & 6'd21
                                | {6{gpr17_recover_table[22]}} & 6'd22
                                | {6{gpr17_recover_table[23]}} & 6'd23
                                | {6{gpr17_recover_table[24]}} & 6'd24
                                | {6{gpr17_recover_table[25]}} & 6'd25
                                | {6{gpr17_recover_table[26]}} & 6'd26
                                | {6{gpr17_recover_table[27]}} & 6'd27
                                | {6{gpr17_recover_table[28]}} & 6'd28
                                | {6{gpr17_recover_table[29]}} & 6'd29
                                | {6{gpr17_recover_table[30]}} & 6'd30
                                | {6{gpr17_recover_table[31]}} & 6'd31
                                | {6{gpr17_recover_table[32]}} & 6'd32
                                | {6{gpr17_recover_table[33]}} & 6'd33
                                | {6{gpr17_recover_table[34]}} & 6'd34
                                | {6{gpr17_recover_table[35]}} & 6'd35
                                | {6{gpr17_recover_table[36]}} & 6'd36
                                | {6{gpr17_recover_table[37]}} & 6'd37
                                | {6{gpr17_recover_table[38]}} & 6'd38
                                | {6{gpr17_recover_table[39]}} & 6'd39
                                | {6{gpr17_recover_table[40]}} & 6'd40
                                | {6{gpr17_recover_table[41]}} & 6'd41
                                | {6{gpr17_recover_table[42]}} & 6'd42
                                | {6{gpr17_recover_table[43]}} & 6'd43
                                | {6{gpr17_recover_table[44]}} & 6'd44
                                | {6{gpr17_recover_table[45]}} & 6'd45
                                | {6{gpr17_recover_table[46]}} & 6'd46
                                | {6{gpr17_recover_table[47]}} & 6'd47
                                | {6{gpr17_recover_table[48]}} & 6'd48
                                | {6{gpr17_recover_table[49]}} & 6'd49
                                | {6{gpr17_recover_table[50]}} & 6'd50
                                | {6{gpr17_recover_table[51]}} & 6'd51
                                | {6{gpr17_recover_table[52]}} & 6'd52
                                | {6{gpr17_recover_table[53]}} & 6'd53
                                | {6{gpr17_recover_table[54]}} & 6'd54
                                | {6{gpr17_recover_table[55]}} & 6'd55
                                | {6{gpr17_recover_table[56]}} & 6'd56
                                | {6{gpr17_recover_table[57]}} & 6'd57
                                | {6{gpr17_recover_table[58]}} & 6'd58
                                | {6{gpr17_recover_table[59]}} & 6'd59
                                | {6{gpr17_recover_table[60]}} & 6'd60
                                | {6{gpr17_recover_table[61]}} & 6'd61
                                | {6{gpr17_recover_table[62]}} & 6'd62
                                | {6{gpr17_recover_table[63]}} & 6'd63;
    assign gpr18_recover_mapped = {6{gpr18_recover_table[0]}}  & 6'd0
                                | {6{gpr18_recover_table[1]}}  & 6'd1
                                | {6{gpr18_recover_table[2]}}  & 6'd2
                                | {6{gpr18_recover_table[3]}}  & 6'd3
                                | {6{gpr18_recover_table[4]}}  & 6'd4
                                | {6{gpr18_recover_table[5]}}  & 6'd5
                                | {6{gpr18_recover_table[6]}}  & 6'd6
                                | {6{gpr18_recover_table[7]}}  & 6'd7
                                | {6{gpr18_recover_table[8]}}  & 6'd8
                                | {6{gpr18_recover_table[9]}}  & 6'd9
                                | {6{gpr18_recover_table[10]}} & 6'd10
                                | {6{gpr18_recover_table[11]}} & 6'd11
                                | {6{gpr18_recover_table[12]}} & 6'd12
                                | {6{gpr18_recover_table[13]}} & 6'd13
                                | {6{gpr18_recover_table[14]}} & 6'd14
                                | {6{gpr18_recover_table[15]}} & 6'd15
                                | {6{gpr18_recover_table[16]}} & 6'd16
                                | {6{gpr18_recover_table[17]}} & 6'd17
                                | {6{gpr18_recover_table[18]}} & 6'd18
                                | {6{gpr18_recover_table[19]}} & 6'd19
                                | {6{gpr18_recover_table[20]}} & 6'd20
                                | {6{gpr18_recover_table[21]}} & 6'd21
                                | {6{gpr18_recover_table[22]}} & 6'd22
                                | {6{gpr18_recover_table[23]}} & 6'd23
                                | {6{gpr18_recover_table[24]}} & 6'd24
                                | {6{gpr18_recover_table[25]}} & 6'd25
                                | {6{gpr18_recover_table[26]}} & 6'd26
                                | {6{gpr18_recover_table[27]}} & 6'd27
                                | {6{gpr18_recover_table[28]}} & 6'd28
                                | {6{gpr18_recover_table[29]}} & 6'd29
                                | {6{gpr18_recover_table[30]}} & 6'd30
                                | {6{gpr18_recover_table[31]}} & 6'd31
                                | {6{gpr18_recover_table[32]}} & 6'd32
                                | {6{gpr18_recover_table[33]}} & 6'd33
                                | {6{gpr18_recover_table[34]}} & 6'd34
                                | {6{gpr18_recover_table[35]}} & 6'd35
                                | {6{gpr18_recover_table[36]}} & 6'd36
                                | {6{gpr18_recover_table[37]}} & 6'd37
                                | {6{gpr18_recover_table[38]}} & 6'd38
                                | {6{gpr18_recover_table[39]}} & 6'd39
                                | {6{gpr18_recover_table[40]}} & 6'd40
                                | {6{gpr18_recover_table[41]}} & 6'd41
                                | {6{gpr18_recover_table[42]}} & 6'd42
                                | {6{gpr18_recover_table[43]}} & 6'd43
                                | {6{gpr18_recover_table[44]}} & 6'd44
                                | {6{gpr18_recover_table[45]}} & 6'd45
                                | {6{gpr18_recover_table[46]}} & 6'd46
                                | {6{gpr18_recover_table[47]}} & 6'd47
                                | {6{gpr18_recover_table[48]}} & 6'd48
                                | {6{gpr18_recover_table[49]}} & 6'd49
                                | {6{gpr18_recover_table[50]}} & 6'd50
                                | {6{gpr18_recover_table[51]}} & 6'd51
                                | {6{gpr18_recover_table[52]}} & 6'd52
                                | {6{gpr18_recover_table[53]}} & 6'd53
                                | {6{gpr18_recover_table[54]}} & 6'd54
                                | {6{gpr18_recover_table[55]}} & 6'd55
                                | {6{gpr18_recover_table[56]}} & 6'd56
                                | {6{gpr18_recover_table[57]}} & 6'd57
                                | {6{gpr18_recover_table[58]}} & 6'd58
                                | {6{gpr18_recover_table[59]}} & 6'd59
                                | {6{gpr18_recover_table[60]}} & 6'd60
                                | {6{gpr18_recover_table[61]}} & 6'd61
                                | {6{gpr18_recover_table[62]}} & 6'd62
                                | {6{gpr18_recover_table[63]}} & 6'd63;
    assign gpr19_recover_mapped = {6{gpr19_recover_table[0]}}  & 6'd0
                                | {6{gpr19_recover_table[1]}}  & 6'd1
                                | {6{gpr19_recover_table[2]}}  & 6'd2
                                | {6{gpr19_recover_table[3]}}  & 6'd3
                                | {6{gpr19_recover_table[4]}}  & 6'd4
                                | {6{gpr19_recover_table[5]}}  & 6'd5
                                | {6{gpr19_recover_table[6]}}  & 6'd6
                                | {6{gpr19_recover_table[7]}}  & 6'd7
                                | {6{gpr19_recover_table[8]}}  & 6'd8
                                | {6{gpr19_recover_table[9]}}  & 6'd9
                                | {6{gpr19_recover_table[10]}} & 6'd10
                                | {6{gpr19_recover_table[11]}} & 6'd11
                                | {6{gpr19_recover_table[12]}} & 6'd12
                                | {6{gpr19_recover_table[13]}} & 6'd13
                                | {6{gpr19_recover_table[14]}} & 6'd14
                                | {6{gpr19_recover_table[15]}} & 6'd15
                                | {6{gpr19_recover_table[16]}} & 6'd16
                                | {6{gpr19_recover_table[17]}} & 6'd17
                                | {6{gpr19_recover_table[18]}} & 6'd18
                                | {6{gpr19_recover_table[19]}} & 6'd19
                                | {6{gpr19_recover_table[20]}} & 6'd20
                                | {6{gpr19_recover_table[21]}} & 6'd21
                                | {6{gpr19_recover_table[22]}} & 6'd22
                                | {6{gpr19_recover_table[23]}} & 6'd23
                                | {6{gpr19_recover_table[24]}} & 6'd24
                                | {6{gpr19_recover_table[25]}} & 6'd25
                                | {6{gpr19_recover_table[26]}} & 6'd26
                                | {6{gpr19_recover_table[27]}} & 6'd27
                                | {6{gpr19_recover_table[28]}} & 6'd28
                                | {6{gpr19_recover_table[29]}} & 6'd29
                                | {6{gpr19_recover_table[30]}} & 6'd30
                                | {6{gpr19_recover_table[31]}} & 6'd31
                                | {6{gpr19_recover_table[32]}} & 6'd32
                                | {6{gpr19_recover_table[33]}} & 6'd33
                                | {6{gpr19_recover_table[34]}} & 6'd34
                                | {6{gpr19_recover_table[35]}} & 6'd35
                                | {6{gpr19_recover_table[36]}} & 6'd36
                                | {6{gpr19_recover_table[37]}} & 6'd37
                                | {6{gpr19_recover_table[38]}} & 6'd38
                                | {6{gpr19_recover_table[39]}} & 6'd39
                                | {6{gpr19_recover_table[40]}} & 6'd40
                                | {6{gpr19_recover_table[41]}} & 6'd41
                                | {6{gpr19_recover_table[42]}} & 6'd42
                                | {6{gpr19_recover_table[43]}} & 6'd43
                                | {6{gpr19_recover_table[44]}} & 6'd44
                                | {6{gpr19_recover_table[45]}} & 6'd45
                                | {6{gpr19_recover_table[46]}} & 6'd46
                                | {6{gpr19_recover_table[47]}} & 6'd47
                                | {6{gpr19_recover_table[48]}} & 6'd48
                                | {6{gpr19_recover_table[49]}} & 6'd49
                                | {6{gpr19_recover_table[50]}} & 6'd50
                                | {6{gpr19_recover_table[51]}} & 6'd51
                                | {6{gpr19_recover_table[52]}} & 6'd52
                                | {6{gpr19_recover_table[53]}} & 6'd53
                                | {6{gpr19_recover_table[54]}} & 6'd54
                                | {6{gpr19_recover_table[55]}} & 6'd55
                                | {6{gpr19_recover_table[56]}} & 6'd56
                                | {6{gpr19_recover_table[57]}} & 6'd57
                                | {6{gpr19_recover_table[58]}} & 6'd58
                                | {6{gpr19_recover_table[59]}} & 6'd59
                                | {6{gpr19_recover_table[60]}} & 6'd60
                                | {6{gpr19_recover_table[61]}} & 6'd61
                                | {6{gpr19_recover_table[62]}} & 6'd62
                                | {6{gpr19_recover_table[63]}} & 6'd63;
    assign gpr20_recover_mapped = {6{gpr20_recover_table[0]}}  & 6'd0
                                | {6{gpr20_recover_table[1]}}  & 6'd1
                                | {6{gpr20_recover_table[2]}}  & 6'd2
                                | {6{gpr20_recover_table[3]}}  & 6'd3
                                | {6{gpr20_recover_table[4]}}  & 6'd4
                                | {6{gpr20_recover_table[5]}}  & 6'd5
                                | {6{gpr20_recover_table[6]}}  & 6'd6
                                | {6{gpr20_recover_table[7]}}  & 6'd7
                                | {6{gpr20_recover_table[8]}}  & 6'd8
                                | {6{gpr20_recover_table[9]}}  & 6'd9
                                | {6{gpr20_recover_table[10]}} & 6'd10
                                | {6{gpr20_recover_table[11]}} & 6'd11
                                | {6{gpr20_recover_table[12]}} & 6'd12
                                | {6{gpr20_recover_table[13]}} & 6'd13
                                | {6{gpr20_recover_table[14]}} & 6'd14
                                | {6{gpr20_recover_table[15]}} & 6'd15
                                | {6{gpr20_recover_table[16]}} & 6'd16
                                | {6{gpr20_recover_table[17]}} & 6'd17
                                | {6{gpr20_recover_table[18]}} & 6'd18
                                | {6{gpr20_recover_table[19]}} & 6'd19
                                | {6{gpr20_recover_table[20]}} & 6'd20
                                | {6{gpr20_recover_table[21]}} & 6'd21
                                | {6{gpr20_recover_table[22]}} & 6'd22
                                | {6{gpr20_recover_table[23]}} & 6'd23
                                | {6{gpr20_recover_table[24]}} & 6'd24
                                | {6{gpr20_recover_table[25]}} & 6'd25
                                | {6{gpr20_recover_table[26]}} & 6'd26
                                | {6{gpr20_recover_table[27]}} & 6'd27
                                | {6{gpr20_recover_table[28]}} & 6'd28
                                | {6{gpr20_recover_table[29]}} & 6'd29
                                | {6{gpr20_recover_table[30]}} & 6'd30
                                | {6{gpr20_recover_table[31]}} & 6'd31
                                | {6{gpr20_recover_table[32]}} & 6'd32
                                | {6{gpr20_recover_table[33]}} & 6'd33
                                | {6{gpr20_recover_table[34]}} & 6'd34
                                | {6{gpr20_recover_table[35]}} & 6'd35
                                | {6{gpr20_recover_table[36]}} & 6'd36
                                | {6{gpr20_recover_table[37]}} & 6'd37
                                | {6{gpr20_recover_table[38]}} & 6'd38
                                | {6{gpr20_recover_table[39]}} & 6'd39
                                | {6{gpr20_recover_table[40]}} & 6'd40
                                | {6{gpr20_recover_table[41]}} & 6'd41
                                | {6{gpr20_recover_table[42]}} & 6'd42
                                | {6{gpr20_recover_table[43]}} & 6'd43
                                | {6{gpr20_recover_table[44]}} & 6'd44
                                | {6{gpr20_recover_table[45]}} & 6'd45
                                | {6{gpr20_recover_table[46]}} & 6'd46
                                | {6{gpr20_recover_table[47]}} & 6'd47
                                | {6{gpr20_recover_table[48]}} & 6'd48
                                | {6{gpr20_recover_table[49]}} & 6'd49
                                | {6{gpr20_recover_table[50]}} & 6'd50
                                | {6{gpr20_recover_table[51]}} & 6'd51
                                | {6{gpr20_recover_table[52]}} & 6'd52
                                | {6{gpr20_recover_table[53]}} & 6'd53
                                | {6{gpr20_recover_table[54]}} & 6'd54
                                | {6{gpr20_recover_table[55]}} & 6'd55
                                | {6{gpr20_recover_table[56]}} & 6'd56
                                | {6{gpr20_recover_table[57]}} & 6'd57
                                | {6{gpr20_recover_table[58]}} & 6'd58
                                | {6{gpr20_recover_table[59]}} & 6'd59
                                | {6{gpr20_recover_table[60]}} & 6'd60
                                | {6{gpr20_recover_table[61]}} & 6'd61
                                | {6{gpr20_recover_table[62]}} & 6'd62
                                | {6{gpr20_recover_table[63]}} & 6'd63;
    assign gpr21_recover_mapped = {6{gpr21_recover_table[0]}}  & 6'd0
                                | {6{gpr21_recover_table[1]}}  & 6'd1
                                | {6{gpr21_recover_table[2]}}  & 6'd2
                                | {6{gpr21_recover_table[3]}}  & 6'd3
                                | {6{gpr21_recover_table[4]}}  & 6'd4
                                | {6{gpr21_recover_table[5]}}  & 6'd5
                                | {6{gpr21_recover_table[6]}}  & 6'd6
                                | {6{gpr21_recover_table[7]}}  & 6'd7
                                | {6{gpr21_recover_table[8]}}  & 6'd8
                                | {6{gpr21_recover_table[9]}}  & 6'd9
                                | {6{gpr21_recover_table[10]}} & 6'd10
                                | {6{gpr21_recover_table[11]}} & 6'd11
                                | {6{gpr21_recover_table[12]}} & 6'd12
                                | {6{gpr21_recover_table[13]}} & 6'd13
                                | {6{gpr21_recover_table[14]}} & 6'd14
                                | {6{gpr21_recover_table[15]}} & 6'd15
                                | {6{gpr21_recover_table[16]}} & 6'd16
                                | {6{gpr21_recover_table[17]}} & 6'd17
                                | {6{gpr21_recover_table[18]}} & 6'd18
                                | {6{gpr21_recover_table[19]}} & 6'd19
                                | {6{gpr21_recover_table[20]}} & 6'd20
                                | {6{gpr21_recover_table[21]}} & 6'd21
                                | {6{gpr21_recover_table[22]}} & 6'd22
                                | {6{gpr21_recover_table[23]}} & 6'd23
                                | {6{gpr21_recover_table[24]}} & 6'd24
                                | {6{gpr21_recover_table[25]}} & 6'd25
                                | {6{gpr21_recover_table[26]}} & 6'd26
                                | {6{gpr21_recover_table[27]}} & 6'd27
                                | {6{gpr21_recover_table[28]}} & 6'd28
                                | {6{gpr21_recover_table[29]}} & 6'd29
                                | {6{gpr21_recover_table[30]}} & 6'd30
                                | {6{gpr21_recover_table[31]}} & 6'd31
                                | {6{gpr21_recover_table[32]}} & 6'd32
                                | {6{gpr21_recover_table[33]}} & 6'd33
                                | {6{gpr21_recover_table[34]}} & 6'd34
                                | {6{gpr21_recover_table[35]}} & 6'd35
                                | {6{gpr21_recover_table[36]}} & 6'd36
                                | {6{gpr21_recover_table[37]}} & 6'd37
                                | {6{gpr21_recover_table[38]}} & 6'd38
                                | {6{gpr21_recover_table[39]}} & 6'd39
                                | {6{gpr21_recover_table[40]}} & 6'd40
                                | {6{gpr21_recover_table[41]}} & 6'd41
                                | {6{gpr21_recover_table[42]}} & 6'd42
                                | {6{gpr21_recover_table[43]}} & 6'd43
                                | {6{gpr21_recover_table[44]}} & 6'd44
                                | {6{gpr21_recover_table[45]}} & 6'd45
                                | {6{gpr21_recover_table[46]}} & 6'd46
                                | {6{gpr21_recover_table[47]}} & 6'd47
                                | {6{gpr21_recover_table[48]}} & 6'd48
                                | {6{gpr21_recover_table[49]}} & 6'd49
                                | {6{gpr21_recover_table[50]}} & 6'd50
                                | {6{gpr21_recover_table[51]}} & 6'd51
                                | {6{gpr21_recover_table[52]}} & 6'd52
                                | {6{gpr21_recover_table[53]}} & 6'd53
                                | {6{gpr21_recover_table[54]}} & 6'd54
                                | {6{gpr21_recover_table[55]}} & 6'd55
                                | {6{gpr21_recover_table[56]}} & 6'd56
                                | {6{gpr21_recover_table[57]}} & 6'd57
                                | {6{gpr21_recover_table[58]}} & 6'd58
                                | {6{gpr21_recover_table[59]}} & 6'd59
                                | {6{gpr21_recover_table[60]}} & 6'd60
                                | {6{gpr21_recover_table[61]}} & 6'd61
                                | {6{gpr21_recover_table[62]}} & 6'd62
                                | {6{gpr21_recover_table[63]}} & 6'd63;
    assign gpr22_recover_mapped = {6{gpr22_recover_table[0]}}  & 6'd0
                                | {6{gpr22_recover_table[1]}}  & 6'd1
                                | {6{gpr22_recover_table[2]}}  & 6'd2
                                | {6{gpr22_recover_table[3]}}  & 6'd3
                                | {6{gpr22_recover_table[4]}}  & 6'd4
                                | {6{gpr22_recover_table[5]}}  & 6'd5
                                | {6{gpr22_recover_table[6]}}  & 6'd6
                                | {6{gpr22_recover_table[7]}}  & 6'd7
                                | {6{gpr22_recover_table[8]}}  & 6'd8
                                | {6{gpr22_recover_table[9]}}  & 6'd9
                                | {6{gpr22_recover_table[10]}} & 6'd10
                                | {6{gpr22_recover_table[11]}} & 6'd11
                                | {6{gpr22_recover_table[12]}} & 6'd12
                                | {6{gpr22_recover_table[13]}} & 6'd13
                                | {6{gpr22_recover_table[14]}} & 6'd14
                                | {6{gpr22_recover_table[15]}} & 6'd15
                                | {6{gpr22_recover_table[16]}} & 6'd16
                                | {6{gpr22_recover_table[17]}} & 6'd17
                                | {6{gpr22_recover_table[18]}} & 6'd18
                                | {6{gpr22_recover_table[19]}} & 6'd19
                                | {6{gpr22_recover_table[20]}} & 6'd20
                                | {6{gpr22_recover_table[21]}} & 6'd21
                                | {6{gpr22_recover_table[22]}} & 6'd22
                                | {6{gpr22_recover_table[23]}} & 6'd23
                                | {6{gpr22_recover_table[24]}} & 6'd24
                                | {6{gpr22_recover_table[25]}} & 6'd25
                                | {6{gpr22_recover_table[26]}} & 6'd26
                                | {6{gpr22_recover_table[27]}} & 6'd27
                                | {6{gpr22_recover_table[28]}} & 6'd28
                                | {6{gpr22_recover_table[29]}} & 6'd29
                                | {6{gpr22_recover_table[30]}} & 6'd30
                                | {6{gpr22_recover_table[31]}} & 6'd31
                                | {6{gpr22_recover_table[32]}} & 6'd32
                                | {6{gpr22_recover_table[33]}} & 6'd33
                                | {6{gpr22_recover_table[34]}} & 6'd34
                                | {6{gpr22_recover_table[35]}} & 6'd35
                                | {6{gpr22_recover_table[36]}} & 6'd36
                                | {6{gpr22_recover_table[37]}} & 6'd37
                                | {6{gpr22_recover_table[38]}} & 6'd38
                                | {6{gpr22_recover_table[39]}} & 6'd39
                                | {6{gpr22_recover_table[40]}} & 6'd40
                                | {6{gpr22_recover_table[41]}} & 6'd41
                                | {6{gpr22_recover_table[42]}} & 6'd42
                                | {6{gpr22_recover_table[43]}} & 6'd43
                                | {6{gpr22_recover_table[44]}} & 6'd44
                                | {6{gpr22_recover_table[45]}} & 6'd45
                                | {6{gpr22_recover_table[46]}} & 6'd46
                                | {6{gpr22_recover_table[47]}} & 6'd47
                                | {6{gpr22_recover_table[48]}} & 6'd48
                                | {6{gpr22_recover_table[49]}} & 6'd49
                                | {6{gpr22_recover_table[50]}} & 6'd50
                                | {6{gpr22_recover_table[51]}} & 6'd51
                                | {6{gpr22_recover_table[52]}} & 6'd52
                                | {6{gpr22_recover_table[53]}} & 6'd53
                                | {6{gpr22_recover_table[54]}} & 6'd54
                                | {6{gpr22_recover_table[55]}} & 6'd55
                                | {6{gpr22_recover_table[56]}} & 6'd56
                                | {6{gpr22_recover_table[57]}} & 6'd57
                                | {6{gpr22_recover_table[58]}} & 6'd58
                                | {6{gpr22_recover_table[59]}} & 6'd59
                                | {6{gpr22_recover_table[60]}} & 6'd60
                                | {6{gpr22_recover_table[61]}} & 6'd61
                                | {6{gpr22_recover_table[62]}} & 6'd62
                                | {6{gpr22_recover_table[63]}} & 6'd63;
    assign gpr23_recover_mapped = {6{gpr23_recover_table[0]}}  & 6'd0
                                | {6{gpr23_recover_table[1]}}  & 6'd1
                                | {6{gpr23_recover_table[2]}}  & 6'd2
                                | {6{gpr23_recover_table[3]}}  & 6'd3
                                | {6{gpr23_recover_table[4]}}  & 6'd4
                                | {6{gpr23_recover_table[5]}}  & 6'd5
                                | {6{gpr23_recover_table[6]}}  & 6'd6
                                | {6{gpr23_recover_table[7]}}  & 6'd7
                                | {6{gpr23_recover_table[8]}}  & 6'd8
                                | {6{gpr23_recover_table[9]}}  & 6'd9
                                | {6{gpr23_recover_table[10]}} & 6'd10
                                | {6{gpr23_recover_table[11]}} & 6'd11
                                | {6{gpr23_recover_table[12]}} & 6'd12
                                | {6{gpr23_recover_table[13]}} & 6'd13
                                | {6{gpr23_recover_table[14]}} & 6'd14
                                | {6{gpr23_recover_table[15]}} & 6'd15
                                | {6{gpr23_recover_table[16]}} & 6'd16
                                | {6{gpr23_recover_table[17]}} & 6'd17
                                | {6{gpr23_recover_table[18]}} & 6'd18
                                | {6{gpr23_recover_table[19]}} & 6'd19
                                | {6{gpr23_recover_table[20]}} & 6'd20
                                | {6{gpr23_recover_table[21]}} & 6'd21
                                | {6{gpr23_recover_table[22]}} & 6'd22
                                | {6{gpr23_recover_table[23]}} & 6'd23
                                | {6{gpr23_recover_table[24]}} & 6'd24
                                | {6{gpr23_recover_table[25]}} & 6'd25
                                | {6{gpr23_recover_table[26]}} & 6'd26
                                | {6{gpr23_recover_table[27]}} & 6'd27
                                | {6{gpr23_recover_table[28]}} & 6'd28
                                | {6{gpr23_recover_table[29]}} & 6'd29
                                | {6{gpr23_recover_table[30]}} & 6'd30
                                | {6{gpr23_recover_table[31]}} & 6'd31
                                | {6{gpr23_recover_table[32]}} & 6'd32
                                | {6{gpr23_recover_table[33]}} & 6'd33
                                | {6{gpr23_recover_table[34]}} & 6'd34
                                | {6{gpr23_recover_table[35]}} & 6'd35
                                | {6{gpr23_recover_table[36]}} & 6'd36
                                | {6{gpr23_recover_table[37]}} & 6'd37
                                | {6{gpr23_recover_table[38]}} & 6'd38
                                | {6{gpr23_recover_table[39]}} & 6'd39
                                | {6{gpr23_recover_table[40]}} & 6'd40
                                | {6{gpr23_recover_table[41]}} & 6'd41
                                | {6{gpr23_recover_table[42]}} & 6'd42
                                | {6{gpr23_recover_table[43]}} & 6'd43
                                | {6{gpr23_recover_table[44]}} & 6'd44
                                | {6{gpr23_recover_table[45]}} & 6'd45
                                | {6{gpr23_recover_table[46]}} & 6'd46
                                | {6{gpr23_recover_table[47]}} & 6'd47
                                | {6{gpr23_recover_table[48]}} & 6'd48
                                | {6{gpr23_recover_table[49]}} & 6'd49
                                | {6{gpr23_recover_table[50]}} & 6'd50
                                | {6{gpr23_recover_table[51]}} & 6'd51
                                | {6{gpr23_recover_table[52]}} & 6'd52
                                | {6{gpr23_recover_table[53]}} & 6'd53
                                | {6{gpr23_recover_table[54]}} & 6'd54
                                | {6{gpr23_recover_table[55]}} & 6'd55
                                | {6{gpr23_recover_table[56]}} & 6'd56
                                | {6{gpr23_recover_table[57]}} & 6'd57
                                | {6{gpr23_recover_table[58]}} & 6'd58
                                | {6{gpr23_recover_table[59]}} & 6'd59
                                | {6{gpr23_recover_table[60]}} & 6'd60
                                | {6{gpr23_recover_table[61]}} & 6'd61
                                | {6{gpr23_recover_table[62]}} & 6'd62
                                | {6{gpr23_recover_table[63]}} & 6'd63;
    assign gpr24_recover_mapped = {6{gpr24_recover_table[0]}}  & 6'd0
                                | {6{gpr24_recover_table[1]}}  & 6'd1
                                | {6{gpr24_recover_table[2]}}  & 6'd2
                                | {6{gpr24_recover_table[3]}}  & 6'd3
                                | {6{gpr24_recover_table[4]}}  & 6'd4
                                | {6{gpr24_recover_table[5]}}  & 6'd5
                                | {6{gpr24_recover_table[6]}}  & 6'd6
                                | {6{gpr24_recover_table[7]}}  & 6'd7
                                | {6{gpr24_recover_table[8]}}  & 6'd8
                                | {6{gpr24_recover_table[9]}}  & 6'd9
                                | {6{gpr24_recover_table[10]}} & 6'd10
                                | {6{gpr24_recover_table[11]}} & 6'd11
                                | {6{gpr24_recover_table[12]}} & 6'd12
                                | {6{gpr24_recover_table[13]}} & 6'd13
                                | {6{gpr24_recover_table[14]}} & 6'd14
                                | {6{gpr24_recover_table[15]}} & 6'd15
                                | {6{gpr24_recover_table[16]}} & 6'd16
                                | {6{gpr24_recover_table[17]}} & 6'd17
                                | {6{gpr24_recover_table[18]}} & 6'd18
                                | {6{gpr24_recover_table[19]}} & 6'd19
                                | {6{gpr24_recover_table[20]}} & 6'd20
                                | {6{gpr24_recover_table[21]}} & 6'd21
                                | {6{gpr24_recover_table[22]}} & 6'd22
                                | {6{gpr24_recover_table[23]}} & 6'd23
                                | {6{gpr24_recover_table[24]}} & 6'd24
                                | {6{gpr24_recover_table[25]}} & 6'd25
                                | {6{gpr24_recover_table[26]}} & 6'd26
                                | {6{gpr24_recover_table[27]}} & 6'd27
                                | {6{gpr24_recover_table[28]}} & 6'd28
                                | {6{gpr24_recover_table[29]}} & 6'd29
                                | {6{gpr24_recover_table[30]}} & 6'd30
                                | {6{gpr24_recover_table[31]}} & 6'd31
                                | {6{gpr24_recover_table[32]}} & 6'd32
                                | {6{gpr24_recover_table[33]}} & 6'd33
                                | {6{gpr24_recover_table[34]}} & 6'd34
                                | {6{gpr24_recover_table[35]}} & 6'd35
                                | {6{gpr24_recover_table[36]}} & 6'd36
                                | {6{gpr24_recover_table[37]}} & 6'd37
                                | {6{gpr24_recover_table[38]}} & 6'd38
                                | {6{gpr24_recover_table[39]}} & 6'd39
                                | {6{gpr24_recover_table[40]}} & 6'd40
                                | {6{gpr24_recover_table[41]}} & 6'd41
                                | {6{gpr24_recover_table[42]}} & 6'd42
                                | {6{gpr24_recover_table[43]}} & 6'd43
                                | {6{gpr24_recover_table[44]}} & 6'd44
                                | {6{gpr24_recover_table[45]}} & 6'd45
                                | {6{gpr24_recover_table[46]}} & 6'd46
                                | {6{gpr24_recover_table[47]}} & 6'd47
                                | {6{gpr24_recover_table[48]}} & 6'd48
                                | {6{gpr24_recover_table[49]}} & 6'd49
                                | {6{gpr24_recover_table[50]}} & 6'd50
                                | {6{gpr24_recover_table[51]}} & 6'd51
                                | {6{gpr24_recover_table[52]}} & 6'd52
                                | {6{gpr24_recover_table[53]}} & 6'd53
                                | {6{gpr24_recover_table[54]}} & 6'd54
                                | {6{gpr24_recover_table[55]}} & 6'd55
                                | {6{gpr24_recover_table[56]}} & 6'd56
                                | {6{gpr24_recover_table[57]}} & 6'd57
                                | {6{gpr24_recover_table[58]}} & 6'd58
                                | {6{gpr24_recover_table[59]}} & 6'd59
                                | {6{gpr24_recover_table[60]}} & 6'd60
                                | {6{gpr24_recover_table[61]}} & 6'd61
                                | {6{gpr24_recover_table[62]}} & 6'd62
                                | {6{gpr24_recover_table[63]}} & 6'd63;
    assign gpr25_recover_mapped = {6{gpr25_recover_table[0]}}  & 6'd0
                                | {6{gpr25_recover_table[1]}}  & 6'd1
                                | {6{gpr25_recover_table[2]}}  & 6'd2
                                | {6{gpr25_recover_table[3]}}  & 6'd3
                                | {6{gpr25_recover_table[4]}}  & 6'd4
                                | {6{gpr25_recover_table[5]}}  & 6'd5
                                | {6{gpr25_recover_table[6]}}  & 6'd6
                                | {6{gpr25_recover_table[7]}}  & 6'd7
                                | {6{gpr25_recover_table[8]}}  & 6'd8
                                | {6{gpr25_recover_table[9]}}  & 6'd9
                                | {6{gpr25_recover_table[10]}} & 6'd10
                                | {6{gpr25_recover_table[11]}} & 6'd11
                                | {6{gpr25_recover_table[12]}} & 6'd12
                                | {6{gpr25_recover_table[13]}} & 6'd13
                                | {6{gpr25_recover_table[14]}} & 6'd14
                                | {6{gpr25_recover_table[15]}} & 6'd15
                                | {6{gpr25_recover_table[16]}} & 6'd16
                                | {6{gpr25_recover_table[17]}} & 6'd17
                                | {6{gpr25_recover_table[18]}} & 6'd18
                                | {6{gpr25_recover_table[19]}} & 6'd19
                                | {6{gpr25_recover_table[20]}} & 6'd20
                                | {6{gpr25_recover_table[21]}} & 6'd21
                                | {6{gpr25_recover_table[22]}} & 6'd22
                                | {6{gpr25_recover_table[23]}} & 6'd23
                                | {6{gpr25_recover_table[24]}} & 6'd24
                                | {6{gpr25_recover_table[25]}} & 6'd25
                                | {6{gpr25_recover_table[26]}} & 6'd26
                                | {6{gpr25_recover_table[27]}} & 6'd27
                                | {6{gpr25_recover_table[28]}} & 6'd28
                                | {6{gpr25_recover_table[29]}} & 6'd29
                                | {6{gpr25_recover_table[30]}} & 6'd30
                                | {6{gpr25_recover_table[31]}} & 6'd31
                                | {6{gpr25_recover_table[32]}} & 6'd32
                                | {6{gpr25_recover_table[33]}} & 6'd33
                                | {6{gpr25_recover_table[34]}} & 6'd34
                                | {6{gpr25_recover_table[35]}} & 6'd35
                                | {6{gpr25_recover_table[36]}} & 6'd36
                                | {6{gpr25_recover_table[37]}} & 6'd37
                                | {6{gpr25_recover_table[38]}} & 6'd38
                                | {6{gpr25_recover_table[39]}} & 6'd39
                                | {6{gpr25_recover_table[40]}} & 6'd40
                                | {6{gpr25_recover_table[41]}} & 6'd41
                                | {6{gpr25_recover_table[42]}} & 6'd42
                                | {6{gpr25_recover_table[43]}} & 6'd43
                                | {6{gpr25_recover_table[44]}} & 6'd44
                                | {6{gpr25_recover_table[45]}} & 6'd45
                                | {6{gpr25_recover_table[46]}} & 6'd46
                                | {6{gpr25_recover_table[47]}} & 6'd47
                                | {6{gpr25_recover_table[48]}} & 6'd48
                                | {6{gpr25_recover_table[49]}} & 6'd49
                                | {6{gpr25_recover_table[50]}} & 6'd50
                                | {6{gpr25_recover_table[51]}} & 6'd51
                                | {6{gpr25_recover_table[52]}} & 6'd52
                                | {6{gpr25_recover_table[53]}} & 6'd53
                                | {6{gpr25_recover_table[54]}} & 6'd54
                                | {6{gpr25_recover_table[55]}} & 6'd55
                                | {6{gpr25_recover_table[56]}} & 6'd56
                                | {6{gpr25_recover_table[57]}} & 6'd57
                                | {6{gpr25_recover_table[58]}} & 6'd58
                                | {6{gpr25_recover_table[59]}} & 6'd59
                                | {6{gpr25_recover_table[60]}} & 6'd60
                                | {6{gpr25_recover_table[61]}} & 6'd61
                                | {6{gpr25_recover_table[62]}} & 6'd62
                                | {6{gpr25_recover_table[63]}} & 6'd63;
    assign gpr26_recover_mapped = {6{gpr26_recover_table[0]}}  & 6'd0
                                | {6{gpr26_recover_table[1]}}  & 6'd1
                                | {6{gpr26_recover_table[2]}}  & 6'd2
                                | {6{gpr26_recover_table[3]}}  & 6'd3
                                | {6{gpr26_recover_table[4]}}  & 6'd4
                                | {6{gpr26_recover_table[5]}}  & 6'd5
                                | {6{gpr26_recover_table[6]}}  & 6'd6
                                | {6{gpr26_recover_table[7]}}  & 6'd7
                                | {6{gpr26_recover_table[8]}}  & 6'd8
                                | {6{gpr26_recover_table[9]}}  & 6'd9
                                | {6{gpr26_recover_table[10]}} & 6'd10
                                | {6{gpr26_recover_table[11]}} & 6'd11
                                | {6{gpr26_recover_table[12]}} & 6'd12
                                | {6{gpr26_recover_table[13]}} & 6'd13
                                | {6{gpr26_recover_table[14]}} & 6'd14
                                | {6{gpr26_recover_table[15]}} & 6'd15
                                | {6{gpr26_recover_table[16]}} & 6'd16
                                | {6{gpr26_recover_table[17]}} & 6'd17
                                | {6{gpr26_recover_table[18]}} & 6'd18
                                | {6{gpr26_recover_table[19]}} & 6'd19
                                | {6{gpr26_recover_table[20]}} & 6'd20
                                | {6{gpr26_recover_table[21]}} & 6'd21
                                | {6{gpr26_recover_table[22]}} & 6'd22
                                | {6{gpr26_recover_table[23]}} & 6'd23
                                | {6{gpr26_recover_table[24]}} & 6'd24
                                | {6{gpr26_recover_table[25]}} & 6'd25
                                | {6{gpr26_recover_table[26]}} & 6'd26
                                | {6{gpr26_recover_table[27]}} & 6'd27
                                | {6{gpr26_recover_table[28]}} & 6'd28
                                | {6{gpr26_recover_table[29]}} & 6'd29
                                | {6{gpr26_recover_table[30]}} & 6'd30
                                | {6{gpr26_recover_table[31]}} & 6'd31
                                | {6{gpr26_recover_table[32]}} & 6'd32
                                | {6{gpr26_recover_table[33]}} & 6'd33
                                | {6{gpr26_recover_table[34]}} & 6'd34
                                | {6{gpr26_recover_table[35]}} & 6'd35
                                | {6{gpr26_recover_table[36]}} & 6'd36
                                | {6{gpr26_recover_table[37]}} & 6'd37
                                | {6{gpr26_recover_table[38]}} & 6'd38
                                | {6{gpr26_recover_table[39]}} & 6'd39
                                | {6{gpr26_recover_table[40]}} & 6'd40
                                | {6{gpr26_recover_table[41]}} & 6'd41
                                | {6{gpr26_recover_table[42]}} & 6'd42
                                | {6{gpr26_recover_table[43]}} & 6'd43
                                | {6{gpr26_recover_table[44]}} & 6'd44
                                | {6{gpr26_recover_table[45]}} & 6'd45
                                | {6{gpr26_recover_table[46]}} & 6'd46
                                | {6{gpr26_recover_table[47]}} & 6'd47
                                | {6{gpr26_recover_table[48]}} & 6'd48
                                | {6{gpr26_recover_table[49]}} & 6'd49
                                | {6{gpr26_recover_table[50]}} & 6'd50
                                | {6{gpr26_recover_table[51]}} & 6'd51
                                | {6{gpr26_recover_table[52]}} & 6'd52
                                | {6{gpr26_recover_table[53]}} & 6'd53
                                | {6{gpr26_recover_table[54]}} & 6'd54
                                | {6{gpr26_recover_table[55]}} & 6'd55
                                | {6{gpr26_recover_table[56]}} & 6'd56
                                | {6{gpr26_recover_table[57]}} & 6'd57
                                | {6{gpr26_recover_table[58]}} & 6'd58
                                | {6{gpr26_recover_table[59]}} & 6'd59
                                | {6{gpr26_recover_table[60]}} & 6'd60
                                | {6{gpr26_recover_table[61]}} & 6'd61
                                | {6{gpr26_recover_table[62]}} & 6'd62
                                | {6{gpr26_recover_table[63]}} & 6'd63;
    assign gpr27_recover_mapped = {6{gpr27_recover_table[0]}}  & 6'd0
                                | {6{gpr27_recover_table[1]}}  & 6'd1
                                | {6{gpr27_recover_table[2]}}  & 6'd2
                                | {6{gpr27_recover_table[3]}}  & 6'd3
                                | {6{gpr27_recover_table[4]}}  & 6'd4
                                | {6{gpr27_recover_table[5]}}  & 6'd5
                                | {6{gpr27_recover_table[6]}}  & 6'd6
                                | {6{gpr27_recover_table[7]}}  & 6'd7
                                | {6{gpr27_recover_table[8]}}  & 6'd8
                                | {6{gpr27_recover_table[9]}}  & 6'd9
                                | {6{gpr27_recover_table[10]}} & 6'd10
                                | {6{gpr27_recover_table[11]}} & 6'd11
                                | {6{gpr27_recover_table[12]}} & 6'd12
                                | {6{gpr27_recover_table[13]}} & 6'd13
                                | {6{gpr27_recover_table[14]}} & 6'd14
                                | {6{gpr27_recover_table[15]}} & 6'd15
                                | {6{gpr27_recover_table[16]}} & 6'd16
                                | {6{gpr27_recover_table[17]}} & 6'd17
                                | {6{gpr27_recover_table[18]}} & 6'd18
                                | {6{gpr27_recover_table[19]}} & 6'd19
                                | {6{gpr27_recover_table[20]}} & 6'd20
                                | {6{gpr27_recover_table[21]}} & 6'd21
                                | {6{gpr27_recover_table[22]}} & 6'd22
                                | {6{gpr27_recover_table[23]}} & 6'd23
                                | {6{gpr27_recover_table[24]}} & 6'd24
                                | {6{gpr27_recover_table[25]}} & 6'd25
                                | {6{gpr27_recover_table[26]}} & 6'd26
                                | {6{gpr27_recover_table[27]}} & 6'd27
                                | {6{gpr27_recover_table[28]}} & 6'd28
                                | {6{gpr27_recover_table[29]}} & 6'd29
                                | {6{gpr27_recover_table[30]}} & 6'd30
                                | {6{gpr27_recover_table[31]}} & 6'd31
                                | {6{gpr27_recover_table[32]}} & 6'd32
                                | {6{gpr27_recover_table[33]}} & 6'd33
                                | {6{gpr27_recover_table[34]}} & 6'd34
                                | {6{gpr27_recover_table[35]}} & 6'd35
                                | {6{gpr27_recover_table[36]}} & 6'd36
                                | {6{gpr27_recover_table[37]}} & 6'd37
                                | {6{gpr27_recover_table[38]}} & 6'd38
                                | {6{gpr27_recover_table[39]}} & 6'd39
                                | {6{gpr27_recover_table[40]}} & 6'd40
                                | {6{gpr27_recover_table[41]}} & 6'd41
                                | {6{gpr27_recover_table[42]}} & 6'd42
                                | {6{gpr27_recover_table[43]}} & 6'd43
                                | {6{gpr27_recover_table[44]}} & 6'd44
                                | {6{gpr27_recover_table[45]}} & 6'd45
                                | {6{gpr27_recover_table[46]}} & 6'd46
                                | {6{gpr27_recover_table[47]}} & 6'd47
                                | {6{gpr27_recover_table[48]}} & 6'd48
                                | {6{gpr27_recover_table[49]}} & 6'd49
                                | {6{gpr27_recover_table[50]}} & 6'd50
                                | {6{gpr27_recover_table[51]}} & 6'd51
                                | {6{gpr27_recover_table[52]}} & 6'd52
                                | {6{gpr27_recover_table[53]}} & 6'd53
                                | {6{gpr27_recover_table[54]}} & 6'd54
                                | {6{gpr27_recover_table[55]}} & 6'd55
                                | {6{gpr27_recover_table[56]}} & 6'd56
                                | {6{gpr27_recover_table[57]}} & 6'd57
                                | {6{gpr27_recover_table[58]}} & 6'd58
                                | {6{gpr27_recover_table[59]}} & 6'd59
                                | {6{gpr27_recover_table[60]}} & 6'd60
                                | {6{gpr27_recover_table[61]}} & 6'd61
                                | {6{gpr27_recover_table[62]}} & 6'd62
                                | {6{gpr27_recover_table[63]}} & 6'd63;
    assign gpr28_recover_mapped = {6{gpr28_recover_table[0]}}  & 6'd0
                                | {6{gpr28_recover_table[1]}}  & 6'd1
                                | {6{gpr28_recover_table[2]}}  & 6'd2
                                | {6{gpr28_recover_table[3]}}  & 6'd3
                                | {6{gpr28_recover_table[4]}}  & 6'd4
                                | {6{gpr28_recover_table[5]}}  & 6'd5
                                | {6{gpr28_recover_table[6]}}  & 6'd6
                                | {6{gpr28_recover_table[7]}}  & 6'd7
                                | {6{gpr28_recover_table[8]}}  & 6'd8
                                | {6{gpr28_recover_table[9]}}  & 6'd9
                                | {6{gpr28_recover_table[10]}} & 6'd10
                                | {6{gpr28_recover_table[11]}} & 6'd11
                                | {6{gpr28_recover_table[12]}} & 6'd12
                                | {6{gpr28_recover_table[13]}} & 6'd13
                                | {6{gpr28_recover_table[14]}} & 6'd14
                                | {6{gpr28_recover_table[15]}} & 6'd15
                                | {6{gpr28_recover_table[16]}} & 6'd16
                                | {6{gpr28_recover_table[17]}} & 6'd17
                                | {6{gpr28_recover_table[18]}} & 6'd18
                                | {6{gpr28_recover_table[19]}} & 6'd19
                                | {6{gpr28_recover_table[20]}} & 6'd20
                                | {6{gpr28_recover_table[21]}} & 6'd21
                                | {6{gpr28_recover_table[22]}} & 6'd22
                                | {6{gpr28_recover_table[23]}} & 6'd23
                                | {6{gpr28_recover_table[24]}} & 6'd24
                                | {6{gpr28_recover_table[25]}} & 6'd25
                                | {6{gpr28_recover_table[26]}} & 6'd26
                                | {6{gpr28_recover_table[27]}} & 6'd27
                                | {6{gpr28_recover_table[28]}} & 6'd28
                                | {6{gpr28_recover_table[29]}} & 6'd29
                                | {6{gpr28_recover_table[30]}} & 6'd30
                                | {6{gpr28_recover_table[31]}} & 6'd31
                                | {6{gpr28_recover_table[32]}} & 6'd32
                                | {6{gpr28_recover_table[33]}} & 6'd33
                                | {6{gpr28_recover_table[34]}} & 6'd34
                                | {6{gpr28_recover_table[35]}} & 6'd35
                                | {6{gpr28_recover_table[36]}} & 6'd36
                                | {6{gpr28_recover_table[37]}} & 6'd37
                                | {6{gpr28_recover_table[38]}} & 6'd38
                                | {6{gpr28_recover_table[39]}} & 6'd39
                                | {6{gpr28_recover_table[40]}} & 6'd40
                                | {6{gpr28_recover_table[41]}} & 6'd41
                                | {6{gpr28_recover_table[42]}} & 6'd42
                                | {6{gpr28_recover_table[43]}} & 6'd43
                                | {6{gpr28_recover_table[44]}} & 6'd44
                                | {6{gpr28_recover_table[45]}} & 6'd45
                                | {6{gpr28_recover_table[46]}} & 6'd46
                                | {6{gpr28_recover_table[47]}} & 6'd47
                                | {6{gpr28_recover_table[48]}} & 6'd48
                                | {6{gpr28_recover_table[49]}} & 6'd49
                                | {6{gpr28_recover_table[50]}} & 6'd50
                                | {6{gpr28_recover_table[51]}} & 6'd51
                                | {6{gpr28_recover_table[52]}} & 6'd52
                                | {6{gpr28_recover_table[53]}} & 6'd53
                                | {6{gpr28_recover_table[54]}} & 6'd54
                                | {6{gpr28_recover_table[55]}} & 6'd55
                                | {6{gpr28_recover_table[56]}} & 6'd56
                                | {6{gpr28_recover_table[57]}} & 6'd57
                                | {6{gpr28_recover_table[58]}} & 6'd58
                                | {6{gpr28_recover_table[59]}} & 6'd59
                                | {6{gpr28_recover_table[60]}} & 6'd60
                                | {6{gpr28_recover_table[61]}} & 6'd61
                                | {6{gpr28_recover_table[62]}} & 6'd62
                                | {6{gpr28_recover_table[63]}} & 6'd63;
    assign gpr29_recover_mapped = {6{gpr29_recover_table[0]}}  & 6'd0
                                | {6{gpr29_recover_table[1]}}  & 6'd1
                                | {6{gpr29_recover_table[2]}}  & 6'd2
                                | {6{gpr29_recover_table[3]}}  & 6'd3
                                | {6{gpr29_recover_table[4]}}  & 6'd4
                                | {6{gpr29_recover_table[5]}}  & 6'd5
                                | {6{gpr29_recover_table[6]}}  & 6'd6
                                | {6{gpr29_recover_table[7]}}  & 6'd7
                                | {6{gpr29_recover_table[8]}}  & 6'd8
                                | {6{gpr29_recover_table[9]}}  & 6'd9
                                | {6{gpr29_recover_table[10]}} & 6'd10
                                | {6{gpr29_recover_table[11]}} & 6'd11
                                | {6{gpr29_recover_table[12]}} & 6'd12
                                | {6{gpr29_recover_table[13]}} & 6'd13
                                | {6{gpr29_recover_table[14]}} & 6'd14
                                | {6{gpr29_recover_table[15]}} & 6'd15
                                | {6{gpr29_recover_table[16]}} & 6'd16
                                | {6{gpr29_recover_table[17]}} & 6'd17
                                | {6{gpr29_recover_table[18]}} & 6'd18
                                | {6{gpr29_recover_table[19]}} & 6'd19
                                | {6{gpr29_recover_table[20]}} & 6'd20
                                | {6{gpr29_recover_table[21]}} & 6'd21
                                | {6{gpr29_recover_table[22]}} & 6'd22
                                | {6{gpr29_recover_table[23]}} & 6'd23
                                | {6{gpr29_recover_table[24]}} & 6'd24
                                | {6{gpr29_recover_table[25]}} & 6'd25
                                | {6{gpr29_recover_table[26]}} & 6'd26
                                | {6{gpr29_recover_table[27]}} & 6'd27
                                | {6{gpr29_recover_table[28]}} & 6'd28
                                | {6{gpr29_recover_table[29]}} & 6'd29
                                | {6{gpr29_recover_table[30]}} & 6'd30
                                | {6{gpr29_recover_table[31]}} & 6'd31
                                | {6{gpr29_recover_table[32]}} & 6'd32
                                | {6{gpr29_recover_table[33]}} & 6'd33
                                | {6{gpr29_recover_table[34]}} & 6'd34
                                | {6{gpr29_recover_table[35]}} & 6'd35
                                | {6{gpr29_recover_table[36]}} & 6'd36
                                | {6{gpr29_recover_table[37]}} & 6'd37
                                | {6{gpr29_recover_table[38]}} & 6'd38
                                | {6{gpr29_recover_table[39]}} & 6'd39
                                | {6{gpr29_recover_table[40]}} & 6'd40
                                | {6{gpr29_recover_table[41]}} & 6'd41
                                | {6{gpr29_recover_table[42]}} & 6'd42
                                | {6{gpr29_recover_table[43]}} & 6'd43
                                | {6{gpr29_recover_table[44]}} & 6'd44
                                | {6{gpr29_recover_table[45]}} & 6'd45
                                | {6{gpr29_recover_table[46]}} & 6'd46
                                | {6{gpr29_recover_table[47]}} & 6'd47
                                | {6{gpr29_recover_table[48]}} & 6'd48
                                | {6{gpr29_recover_table[49]}} & 6'd49
                                | {6{gpr29_recover_table[50]}} & 6'd50
                                | {6{gpr29_recover_table[51]}} & 6'd51
                                | {6{gpr29_recover_table[52]}} & 6'd52
                                | {6{gpr29_recover_table[53]}} & 6'd53
                                | {6{gpr29_recover_table[54]}} & 6'd54
                                | {6{gpr29_recover_table[55]}} & 6'd55
                                | {6{gpr29_recover_table[56]}} & 6'd56
                                | {6{gpr29_recover_table[57]}} & 6'd57
                                | {6{gpr29_recover_table[58]}} & 6'd58
                                | {6{gpr29_recover_table[59]}} & 6'd59
                                | {6{gpr29_recover_table[60]}} & 6'd60
                                | {6{gpr29_recover_table[61]}} & 6'd61
                                | {6{gpr29_recover_table[62]}} & 6'd62
                                | {6{gpr29_recover_table[63]}} & 6'd63;
    assign gpr30_recover_mapped = {6{gpr30_recover_table[0]}}  & 6'd0
                                | {6{gpr30_recover_table[1]}}  & 6'd1
                                | {6{gpr30_recover_table[2]}}  & 6'd2
                                | {6{gpr30_recover_table[3]}}  & 6'd3
                                | {6{gpr30_recover_table[4]}}  & 6'd4
                                | {6{gpr30_recover_table[5]}}  & 6'd5
                                | {6{gpr30_recover_table[6]}}  & 6'd6
                                | {6{gpr30_recover_table[7]}}  & 6'd7
                                | {6{gpr30_recover_table[8]}}  & 6'd8
                                | {6{gpr30_recover_table[9]}}  & 6'd9
                                | {6{gpr30_recover_table[10]}} & 6'd10
                                | {6{gpr30_recover_table[11]}} & 6'd11
                                | {6{gpr30_recover_table[12]}} & 6'd12
                                | {6{gpr30_recover_table[13]}} & 6'd13
                                | {6{gpr30_recover_table[14]}} & 6'd14
                                | {6{gpr30_recover_table[15]}} & 6'd15
                                | {6{gpr30_recover_table[16]}} & 6'd16
                                | {6{gpr30_recover_table[17]}} & 6'd17
                                | {6{gpr30_recover_table[18]}} & 6'd18
                                | {6{gpr30_recover_table[19]}} & 6'd19
                                | {6{gpr30_recover_table[20]}} & 6'd20
                                | {6{gpr30_recover_table[21]}} & 6'd21
                                | {6{gpr30_recover_table[22]}} & 6'd22
                                | {6{gpr30_recover_table[23]}} & 6'd23
                                | {6{gpr30_recover_table[24]}} & 6'd24
                                | {6{gpr30_recover_table[25]}} & 6'd25
                                | {6{gpr30_recover_table[26]}} & 6'd26
                                | {6{gpr30_recover_table[27]}} & 6'd27
                                | {6{gpr30_recover_table[28]}} & 6'd28
                                | {6{gpr30_recover_table[29]}} & 6'd29
                                | {6{gpr30_recover_table[30]}} & 6'd30
                                | {6{gpr30_recover_table[31]}} & 6'd31
                                | {6{gpr30_recover_table[32]}} & 6'd32
                                | {6{gpr30_recover_table[33]}} & 6'd33
                                | {6{gpr30_recover_table[34]}} & 6'd34
                                | {6{gpr30_recover_table[35]}} & 6'd35
                                | {6{gpr30_recover_table[36]}} & 6'd36
                                | {6{gpr30_recover_table[37]}} & 6'd37
                                | {6{gpr30_recover_table[38]}} & 6'd38
                                | {6{gpr30_recover_table[39]}} & 6'd39
                                | {6{gpr30_recover_table[40]}} & 6'd40
                                | {6{gpr30_recover_table[41]}} & 6'd41
                                | {6{gpr30_recover_table[42]}} & 6'd42
                                | {6{gpr30_recover_table[43]}} & 6'd43
                                | {6{gpr30_recover_table[44]}} & 6'd44
                                | {6{gpr30_recover_table[45]}} & 6'd45
                                | {6{gpr30_recover_table[46]}} & 6'd46
                                | {6{gpr30_recover_table[47]}} & 6'd47
                                | {6{gpr30_recover_table[48]}} & 6'd48
                                | {6{gpr30_recover_table[49]}} & 6'd49
                                | {6{gpr30_recover_table[50]}} & 6'd50
                                | {6{gpr30_recover_table[51]}} & 6'd51
                                | {6{gpr30_recover_table[52]}} & 6'd52
                                | {6{gpr30_recover_table[53]}} & 6'd53
                                | {6{gpr30_recover_table[54]}} & 6'd54
                                | {6{gpr30_recover_table[55]}} & 6'd55
                                | {6{gpr30_recover_table[56]}} & 6'd56
                                | {6{gpr30_recover_table[57]}} & 6'd57
                                | {6{gpr30_recover_table[58]}} & 6'd58
                                | {6{gpr30_recover_table[59]}} & 6'd59
                                | {6{gpr30_recover_table[60]}} & 6'd60
                                | {6{gpr30_recover_table[61]}} & 6'd61
                                | {6{gpr30_recover_table[62]}} & 6'd62
                                | {6{gpr30_recover_table[63]}} & 6'd63;
    assign gpr31_recover_mapped = {6{gpr31_recover_table[0]}}  & 6'd0
                                | {6{gpr31_recover_table[1]}}  & 6'd1
                                | {6{gpr31_recover_table[2]}}  & 6'd2
                                | {6{gpr31_recover_table[3]}}  & 6'd3
                                | {6{gpr31_recover_table[4]}}  & 6'd4
                                | {6{gpr31_recover_table[5]}}  & 6'd5
                                | {6{gpr31_recover_table[6]}}  & 6'd6
                                | {6{gpr31_recover_table[7]}}  & 6'd7
                                | {6{gpr31_recover_table[8]}}  & 6'd8
                                | {6{gpr31_recover_table[9]}}  & 6'd9
                                | {6{gpr31_recover_table[10]}} & 6'd10
                                | {6{gpr31_recover_table[11]}} & 6'd11
                                | {6{gpr31_recover_table[12]}} & 6'd12
                                | {6{gpr31_recover_table[13]}} & 6'd13
                                | {6{gpr31_recover_table[14]}} & 6'd14
                                | {6{gpr31_recover_table[15]}} & 6'd15
                                | {6{gpr31_recover_table[16]}} & 6'd16
                                | {6{gpr31_recover_table[17]}} & 6'd17
                                | {6{gpr31_recover_table[18]}} & 6'd18
                                | {6{gpr31_recover_table[19]}} & 6'd19
                                | {6{gpr31_recover_table[20]}} & 6'd20
                                | {6{gpr31_recover_table[21]}} & 6'd21
                                | {6{gpr31_recover_table[22]}} & 6'd22
                                | {6{gpr31_recover_table[23]}} & 6'd23
                                | {6{gpr31_recover_table[24]}} & 6'd24
                                | {6{gpr31_recover_table[25]}} & 6'd25
                                | {6{gpr31_recover_table[26]}} & 6'd26
                                | {6{gpr31_recover_table[27]}} & 6'd27
                                | {6{gpr31_recover_table[28]}} & 6'd28
                                | {6{gpr31_recover_table[29]}} & 6'd29
                                | {6{gpr31_recover_table[30]}} & 6'd30
                                | {6{gpr31_recover_table[31]}} & 6'd31
                                | {6{gpr31_recover_table[32]}} & 6'd32
                                | {6{gpr31_recover_table[33]}} & 6'd33
                                | {6{gpr31_recover_table[34]}} & 6'd34
                                | {6{gpr31_recover_table[35]}} & 6'd35
                                | {6{gpr31_recover_table[36]}} & 6'd36
                                | {6{gpr31_recover_table[37]}} & 6'd37
                                | {6{gpr31_recover_table[38]}} & 6'd38
                                | {6{gpr31_recover_table[39]}} & 6'd39
                                | {6{gpr31_recover_table[40]}} & 6'd40
                                | {6{gpr31_recover_table[41]}} & 6'd41
                                | {6{gpr31_recover_table[42]}} & 6'd42
                                | {6{gpr31_recover_table[43]}} & 6'd43
                                | {6{gpr31_recover_table[44]}} & 6'd44
                                | {6{gpr31_recover_table[45]}} & 6'd45
                                | {6{gpr31_recover_table[46]}} & 6'd46
                                | {6{gpr31_recover_table[47]}} & 6'd47
                                | {6{gpr31_recover_table[48]}} & 6'd48
                                | {6{gpr31_recover_table[49]}} & 6'd49
                                | {6{gpr31_recover_table[50]}} & 6'd50
                                | {6{gpr31_recover_table[51]}} & 6'd51
                                | {6{gpr31_recover_table[52]}} & 6'd52
                                | {6{gpr31_recover_table[53]}} & 6'd53
                                | {6{gpr31_recover_table[54]}} & 6'd54
                                | {6{gpr31_recover_table[55]}} & 6'd55
                                | {6{gpr31_recover_table[56]}} & 6'd56
                                | {6{gpr31_recover_table[57]}} & 6'd57
                                | {6{gpr31_recover_table[58]}} & 6'd58
                                | {6{gpr31_recover_table[59]}} & 6'd59
                                | {6{gpr31_recover_table[60]}} & 6'd60
                                | {6{gpr31_recover_table[61]}} & 6'd61
                                | {6{gpr31_recover_table[62]}} & 6'd62
                                | {6{gpr31_recover_table[63]}} & 6'd63;

    assign rtu_idu_ir_recover_table = {gpr31_recover_mapped, gpr30_recover_mapped, gpr29_recover_mapped, gpr28_recover_mapped,
                                       gpr27_recover_mapped, gpr26_recover_mapped, gpr25_recover_mapped, gpr24_recover_mapped,
                                       gpr23_recover_mapped, gpr22_recover_mapped, gpr21_recover_mapped, gpr20_recover_mapped,
                                       gpr19_recover_mapped, gpr18_recover_mapped, gpr17_recover_mapped, gpr16_recover_mapped,
                                       gpr15_recover_mapped, gpr14_recover_mapped, gpr13_recover_mapped, gpr12_recover_mapped,
                                       gpr11_recover_mapped, gpr10_recover_mapped, gpr9_recover_mapped,  gpr8_recover_mapped ,
                                       gpr7_recover_mapped,  gpr6_recover_mapped,  gpr5_recover_mapped,  gpr4_recover_mapped ,
                                       gpr3_recover_mapped,  gpr2_recover_mapped,  gpr1_recover_mapped,  gpr0_recover_mapped};

    /*
     * alloc 信号生成
     *
     * 当 idu ir 需要有 alloc 状态下的寄存器，或者上一周期后没有可用的 alloc 态寄存器（reset 或 flush 后）才可以更新
     */
    assign alloc_preg_invalid = idu_rtu_pst_pdst_req_vld || !alloc_preg_vld;
    assign pre_alloc_vld = |preg_pre_alloc_vld[63:0];

    always @(posedge clk or negedge rst_clk)
    begin
        if (!rst_clk) begin
            alloc_preg_vld <= 1'b0;
            alloc_preg     <= 6'b0;
        end
        else if (rtu_global_flush) begin
            alloc_preg_vld <= 1'b0;
            alloc_preg     <= 6'b0;
        end
        else if (alloc_preg_invalid) begin
            alloc_preg_vld <= pre_alloc_vld;
            alloc_preg     <= pre_alloc_preg;
        end
        else begin
            alloc_preg_vld <= alloc_preg_vld;
            alloc_preg     <= pre_alloc_preg;
        end
    end
endmodule
