module idu_rf_pregfile (
    clk,
    rst_clk,
    idu_idu_rf_x_pipe0_psrc1_vld,
    idu_idu_rf_x_pipe0_psrc1,
    idu_idu_rf_x_pipe0_psrc2_vld,
    idu_idu_rf_x_pipe0_psrc2,
    idu_idu_rf_x_pipe1_psrc1_vld,
    idu_idu_rf_x_pipe1_psrc1,
    idu_idu_rf_x_pipe1_psrc2_vld,
    idu_idu_rf_x_pipe1_psrc2,
    idu_idu_rf_x_pipe2_psrc1_vld,
    idu_idu_rf_x_pipe2_psrc1,
    idu_idu_rf_x_pipe2_psrc2_vld,
    idu_idu_rf_x_pipe2_psrc2,
    idu_idu_rf_x_pipe3_psrc1_vld,
    idu_idu_rf_x_pipe3_psrc1,
    idu_idu_rf_x_pipe3_psrc2_vld,
    idu_idu_rf_x_pipe3_psrc2,
    idu_idu_rf_x_pipe4_psrc1_vld,
    idu_idu_rf_x_pipe4_psrc1,
    exu_idu_rf_alu_wb_vld,
    exu_idu_rf_alu_wb_preg,
    exu_idu_rf_alu_wb_data,
    exu_idu_rf_mxu_wb_vld,
    exu_idu_rf_mxu_wb_preg,
    exu_idu_rf_mxu_wb_data,
    exu_idu_rf_div_wb_vld,
    exu_idu_rf_div_wb_preg,
    exu_idu_rf_div_wb_data,
    exu_idu_rf_bju_wb_vld,
    exu_idu_rf_bju_wb_preg,
    exu_idu_rf_bju_wb_data,
    exu_idu_rf_lsu_wb_vld,
    exu_idu_rf_lsu_wb_preg,
    exu_idu_rf_lsu_wb_data,
    idu_idu_rf_x_pipe0_psrc1_value,
    idu_idu_rf_x_pipe0_psrc2_value,
    idu_idu_rf_x_pipe1_psrc1_value,
    idu_idu_rf_x_pipe1_psrc2_value,
    idu_idu_rf_x_pipe2_psrc1_value,
    idu_idu_rf_x_pipe2_psrc2_value,
    idu_idu_rf_x_pipe3_psrc1_value,
    idu_idu_rf_x_pipe3_psrc2_value,
    idu_idu_rf_x_pipe4_psrc1_value,
    idu_rtu_pst_wb_vld
);
    // &Ports;
    input         clk;
    input         rst_clk;
    input         idu_idu_rf_x_pipe0_psrc1_vld;
    input  [5 :0] idu_idu_rf_x_pipe0_psrc1;
    input         idu_idu_rf_x_pipe0_psrc2_vld;
    input  [5 :0] idu_idu_rf_x_pipe0_psrc2;
    input         idu_idu_rf_x_pipe1_psrc1_vld;
    input  [5 :0] idu_idu_rf_x_pipe1_psrc1;
    input         idu_idu_rf_x_pipe1_psrc2_vld;
    input  [5 :0] idu_idu_rf_x_pipe1_psrc2;
    input         idu_idu_rf_x_pipe2_psrc1_vld;
    input  [5 :0] idu_idu_rf_x_pipe2_psrc1;
    input         idu_idu_rf_x_pipe2_psrc2_vld;
    input  [5 :0] idu_idu_rf_x_pipe2_psrc2;
    input         idu_idu_rf_x_pipe3_psrc1_vld;
    input  [5 :0] idu_idu_rf_x_pipe3_psrc1;
    input         idu_idu_rf_x_pipe3_psrc2_vld;
    input  [5 :0] idu_idu_rf_x_pipe3_psrc2;
    input         idu_idu_rf_x_pipe4_psrc1_vld;
    input  [5 :0] idu_idu_rf_x_pipe4_psrc1;
    input         exu_idu_rf_alu_wb_vld;
    input  [5 :0] exu_idu_rf_alu_wb_preg;
    input  [63:0] exu_idu_rf_alu_wb_data;
    input         exu_idu_rf_mxu_wb_vld;
    input  [5 :0] exu_idu_rf_mxu_wb_preg;
    input  [63:0] exu_idu_rf_mxu_wb_data;
    input         exu_idu_rf_div_wb_vld;
    input  [5 :0] exu_idu_rf_div_wb_preg;
    input  [63:0] exu_idu_rf_div_wb_data;
    input         exu_idu_rf_bju_wb_vld;
    input  [5 :0] exu_idu_rf_bju_wb_preg;
    input  [63:0] exu_idu_rf_bju_wb_data;
    input         exu_idu_rf_lsu_wb_vld;
    input  [5 :0] exu_idu_rf_lsu_wb_preg;
    input  [63:0] exu_idu_rf_lsu_wb_data;
    output [63:0] idu_idu_rf_x_pipe0_psrc1_value;
    output [63:0] idu_idu_rf_x_pipe0_psrc2_value;
    output [63:0] idu_idu_rf_x_pipe1_psrc1_value;
    output [63:0] idu_idu_rf_x_pipe1_psrc2_value;
    output [63:0] idu_idu_rf_x_pipe2_psrc1_value;
    output [63:0] idu_idu_rf_x_pipe2_psrc2_value;
    output [63:0] idu_idu_rf_x_pipe3_psrc1_value;
    output [63:0] idu_idu_rf_x_pipe3_psrc2_value;
    output [63:0] idu_idu_rf_x_pipe4_psrc1_value;
    output [63:0] idu_rtu_pst_wb_vld;

    // &Regs;

    // &Wires;
    wire        clk;
    wire        rst_clk;
    wire        idu_idu_rf_x_pipe0_psrc1_vld;
    wire [5 :0] idu_idu_rf_x_pipe0_psrc1;
    wire        idu_idu_rf_x_pipe0_psrc2_vld;
    wire [5 :0] idu_idu_rf_x_pipe0_psrc2;
    wire        idu_idu_rf_x_pipe1_psrc1_vld;
    wire [5 :0] idu_idu_rf_x_pipe1_psrc1;
    wire        idu_idu_rf_x_pipe1_psrc2_vld;
    wire [5 :0] idu_idu_rf_x_pipe1_psrc2;
    wire        idu_idu_rf_x_pipe2_psrc1_vld;
    wire [5 :0] idu_idu_rf_x_pipe2_psrc1;
    wire        idu_idu_rf_x_pipe2_psrc2_vld;
    wire [5 :0] idu_idu_rf_x_pipe2_psrc2;
    wire        idu_idu_rf_x_pipe3_psrc1_vld;
    wire [5 :0] idu_idu_rf_x_pipe3_psrc1;
    wire        idu_idu_rf_x_pipe3_psrc2_vld;
    wire [5 :0] idu_idu_rf_x_pipe3_psrc2;
    wire        idu_idu_rf_x_pipe4_psrc1_vld;
    wire [5 :0] idu_idu_rf_x_pipe4_psrc1;
    wire        exu_idu_rf_alu_wb_vld;
    wire [5 :0] exu_idu_rf_alu_wb_preg;
    wire [63:0] exu_idu_rf_alu_wb_data;
    wire        exu_idu_rf_mxu_wb_vld;
    wire [5 :0] exu_idu_rf_mxu_wb_preg;
    wire [63:0] exu_idu_rf_mxu_wb_data;
    wire        exu_idu_rf_div_wb_vld;
    wire [5 :0] exu_idu_rf_div_wb_preg;
    wire [63:0] exu_idu_rf_div_wb_data;
    wire        exu_idu_rf_bju_wb_vld;
    wire [5 :0] exu_idu_rf_bju_wb_preg;
    wire [63:0] exu_idu_rf_bju_wb_data;
    wire        exu_idu_rf_lsu_wb_vld;
    wire [5 :0] exu_idu_rf_lsu_wb_preg;
    wire [63:0] exu_idu_rf_lsu_wb_data;
    wire [63:0] idu_idu_rf_x_pipe0_psrc1_value;
    wire [63:0] idu_idu_rf_x_pipe0_psrc2_value;
    wire [63:0] idu_idu_rf_x_pipe1_psrc1_value;
    wire [63:0] idu_idu_rf_x_pipe1_psrc2_value;
    wire [63:0] idu_idu_rf_x_pipe2_psrc1_value;
    wire [63:0] idu_idu_rf_x_pipe2_psrc2_value;
    wire [63:0] idu_idu_rf_x_pipe3_psrc1_value;
    wire [63:0] idu_idu_rf_x_pipe3_psrc2_value;
    wire [63:0] idu_idu_rf_x_pipe4_psrc1_value;

    wire [63:0] data0;
    wire [63:0] data1;
    wire [63:0] data2;
    wire [63:0] data3;
    wire [63:0] data4;
    wire [63:0] data5;
    wire [63:0] data6;
    wire [63:0] data7;
    wire [63:0] data8;
    wire [63:0] data9;
    wire [63:0] data10;
    wire [63:0] data11;
    wire [63:0] data12;
    wire [63:0] data13;
    wire [63:0] data14;
    wire [63:0] data15;
    wire [63:0] data16;
    wire [63:0] data17;
    wire [63:0] data18;
    wire [63:0] data19;
    wire [63:0] data20;
    wire [63:0] data21;
    wire [63:0] data22;
    wire [63:0] data23;
    wire [63:0] data24;
    wire [63:0] data25;
    wire [63:0] data26;
    wire [63:0] data27;
    wire [63:0] data28;
    wire [63:0] data29;
    wire [63:0] data30;
    wire [63:0] data31;
    wire [63:0] data32;
    wire [63:0] data33;
    wire [63:0] data34;
    wire [63:0] data35;
    wire [63:0] data36;
    wire [63:0] data37;
    wire [63:0] data38;
    wire [63:0] data39;
    wire [63:0] data40;
    wire [63:0] data41;
    wire [63:0] data42;
    wire [63:0] data43;
    wire [63:0] data44;
    wire [63:0] data45;
    wire [63:0] data46;
    wire [63:0] data47;
    wire [63:0] data48;
    wire [63:0] data49;
    wire [63:0] data50;
    wire [63:0] data51;
    wire [63:0] data52;
    wire [63:0] data53;
    wire [63:0] data54;
    wire [63:0] data55;
    wire [63:0] data56;
    wire [63:0] data57;
    wire [63:0] data58;
    wire [63:0] data59;
    wire [63:0] data60;
    wire [63:0] data61;
    wire [63:0] data62;
    wire [63:0] data63;
    wire [63:0] pipe0_psrc1_decode;
    wire [63:0] pipe0_psrc2_decode;
    wire [63:0] pipe1_psrc1_decode;
    wire [63:0] pipe1_psrc2_decode;
    wire [63:0] pipe2_psrc1_decode;
    wire [63:0] pipe2_psrc2_decode;
    wire [63:0] pipe3_psrc1_decode;
    wire [63:0] pipe3_psrc2_decode;
    wire [63:0] pipe4_psrc1_decode;
    wire [63:0] alu_wb_en;
    wire [63:0] mxu_wb_en;
    wire [63:0] div_wb_en;
    wire [63:0] bju_wb_en;
    wire [63:0] lsu_wb_en;
    wire [63:0] write_en;
    wire [63:0] write_data0;
    wire [63:0] write_data1;
    wire [63:0] write_data2;
    wire [63:0] write_data3;
    wire [63:0] write_data4;
    wire [63:0] write_data5;
    wire [63:0] write_data6;
    wire [63:0] write_data7;
    wire [63:0] write_data8;
    wire [63:0] write_data9;
    wire [63:0] write_data10;
    wire [63:0] write_data11;
    wire [63:0] write_data12;
    wire [63:0] write_data13;
    wire [63:0] write_data14;
    wire [63:0] write_data15;
    wire [63:0] write_data16;
    wire [63:0] write_data17;
    wire [63:0] write_data18;
    wire [63:0] write_data19;
    wire [63:0] write_data20;
    wire [63:0] write_data21;
    wire [63:0] write_data22;
    wire [63:0] write_data23;
    wire [63:0] write_data24;
    wire [63:0] write_data25;
    wire [63:0] write_data26;
    wire [63:0] write_data27;
    wire [63:0] write_data28;
    wire [63:0] write_data29;
    wire [63:0] write_data30;
    wire [63:0] write_data31;
    wire [63:0] write_data32;
    wire [63:0] write_data33;
    wire [63:0] write_data34;
    wire [63:0] write_data35;
    wire [63:0] write_data36;
    wire [63:0] write_data37;
    wire [63:0] write_data38;
    wire [63:0] write_data39;
    wire [63:0] write_data40;
    wire [63:0] write_data41;
    wire [63:0] write_data42;
    wire [63:0] write_data43;
    wire [63:0] write_data44;
    wire [63:0] write_data45;
    wire [63:0] write_data46;
    wire [63:0] write_data47;
    wire [63:0] write_data48;
    wire [63:0] write_data49;
    wire [63:0] write_data50;
    wire [63:0] write_data51;
    wire [63:0] write_data52;
    wire [63:0] write_data53;
    wire [63:0] write_data54;
    wire [63:0] write_data55;
    wire [63:0] write_data56;
    wire [63:0] write_data57;
    wire [63:0] write_data58;
    wire [63:0] write_data59;
    wire [63:0] write_data60;
    wire [63:0] write_data61;
    wire [63:0] write_data62;
    wire [63:0] write_data63;
    wire [63:0] idu_rtu_pst_wb_vld;

    assign data0 = 0;
    assign idu_rtu_pst_wb_vld[0] = 0;

    idu_rf_preg idu_rf_preg1(
        .clk        	( clk                    ),
        .rst_clk    	( rst_clk                ),
        .write_en   	( write_en[1]            ),
        .write_data 	( write_data1            ),
        .data       	( data1                  ),
        .wb_vld     	( idu_rtu_pst_wb_vld[1]  )
    );

    idu_rf_preg idu_rf_preg2(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[2]            ),
        .write_data     ( write_data2            ),
        .data           ( data2                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[2]  )
    );

    idu_rf_preg idu_rf_preg3(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[3]            ),
        .write_data     ( write_data3            ),
        .data           ( data3                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[3]  )
    );

    idu_rf_preg idu_rf_preg4(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[4]            ),
        .write_data     ( write_data4            ),
        .data           ( data4                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[4]  )
    );

    idu_rf_preg idu_rf_preg5(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[5]            ),
        .write_data     ( write_data5            ),
        .data           ( data5                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[5]  )
    );

    idu_rf_preg idu_rf_preg6(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[6]            ),
        .write_data     ( write_data6            ),
        .data           ( data6                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[6]  )
    );

    idu_rf_preg idu_rf_preg7(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[7]            ),
        .write_data     ( write_data7            ),
        .data           ( data7                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[7]  )
    );

    idu_rf_preg idu_rf_preg8(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[8]            ),
        .write_data     ( write_data8            ),
        .data           ( data8                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[8]  )
    );

    idu_rf_preg idu_rf_preg9(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[9]            ),
        .write_data     ( write_data9            ),
        .data           ( data9                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[9]  )
    );

    idu_rf_preg idu_rf_preg10(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[10]            ),
        .write_data     ( write_data10            ),
        .data           ( data10                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[10]  )
    );

    idu_rf_preg idu_rf_preg11(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[11]            ),
        .write_data     ( write_data11            ),
        .data           ( data11                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[11]  )
    );

    idu_rf_preg idu_rf_preg12(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[12]            ),
        .write_data     ( write_data12            ),
        .data           ( data12                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[12]  )
    );

    idu_rf_preg idu_rf_preg13(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[13]            ),
        .write_data     ( write_data13            ),
        .data           ( data13                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[13]  )
    );

    idu_rf_preg idu_rf_preg14(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[14]            ),
        .write_data     ( write_data14            ),
        .data           ( data14                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[14]  )
    );

    idu_rf_preg idu_rf_preg15(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[15]            ),
        .write_data     ( write_data15            ),
        .data           ( data15                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[15]  )
    );

    idu_rf_preg idu_rf_preg16(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[16]            ),
        .write_data     ( write_data16            ),
        .data           ( data16                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[16]  )
    );

    idu_rf_preg idu_rf_preg17(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[17]            ),
        .write_data     ( write_data17            ),
        .data           ( data17                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[17]  )
    );

    idu_rf_preg idu_rf_preg18(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[18]            ),
        .write_data     ( write_data18            ),
        .data           ( data18                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[18]  )
    );

    idu_rf_preg idu_rf_preg19(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[19]            ),
        .write_data     ( write_data19            ),
        .data           ( data19                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[19]  )
    );

    idu_rf_preg idu_rf_preg20(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[20]            ),
        .write_data     ( write_data20            ),
        .data           ( data20                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[20]  )
    );

    idu_rf_preg idu_rf_preg21(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[21]            ),
        .write_data     ( write_data21            ),
        .data           ( data21                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[21]  )
    );

    idu_rf_preg idu_rf_preg22(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[22]            ),
        .write_data     ( write_data22            ),
        .data           ( data22                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[22]  )
    );

    idu_rf_preg idu_rf_preg23(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[23]            ),
        .write_data     ( write_data23            ),
        .data           ( data23                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[23]  )
    );

    idu_rf_preg idu_rf_preg24(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[24]            ),
        .write_data     ( write_data24            ),
        .data           ( data24                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[24]  )
    );

    idu_rf_preg idu_rf_preg25(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[25]            ),
        .write_data     ( write_data25            ),
        .data           ( data25                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[25]  )
    );

    idu_rf_preg idu_rf_preg26(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[26]            ),
        .write_data     ( write_data26            ),
        .data           ( data26                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[26]  )
    );

    idu_rf_preg idu_rf_preg27(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[27]            ),
        .write_data     ( write_data27            ),
        .data           ( data27                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[27]  )
    );

    idu_rf_preg idu_rf_preg28(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[28]            ),
        .write_data     ( write_data28            ),
        .data           ( data28                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[28]  )
    );

    idu_rf_preg idu_rf_preg29(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[29]            ),
        .write_data     ( write_data29            ),
        .data           ( data29                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[29]  )
    );

    idu_rf_preg idu_rf_preg30(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[30]            ),
        .write_data     ( write_data30            ),
        .data           ( data30                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[30]  )
    );

    idu_rf_preg idu_rf_preg31(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[31]            ),
        .write_data     ( write_data31            ),
        .data           ( data31                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[31]  )
    );

    idu_rf_preg idu_rf_preg32(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[32]            ),
        .write_data     ( write_data32            ),
        .data           ( data32                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[32]  )
    );

    idu_rf_preg idu_rf_preg33(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[33]            ),
        .write_data     ( write_data33            ),
        .data           ( data33                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[33]  )
    );

    idu_rf_preg idu_rf_preg34(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[34]            ),
        .write_data     ( write_data34            ),
        .data           ( data34                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[34]  )
    );

    idu_rf_preg idu_rf_preg35(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[35]            ),
        .write_data     ( write_data35            ),
        .data           ( data35                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[35]  )
    );

    idu_rf_preg idu_rf_preg36(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[36]            ),
        .write_data     ( write_data36            ),
        .data           ( data36                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[36]  )
    );

    idu_rf_preg idu_rf_preg37(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[37]            ),
        .write_data     ( write_data37            ),
        .data           ( data37                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[37]  )
    );

    idu_rf_preg idu_rf_preg38(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[38]            ),
        .write_data     ( write_data38            ),
        .data           ( data38                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[38]  )
    );

    idu_rf_preg idu_rf_preg39(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[39]            ),
        .write_data     ( write_data39            ),
        .data           ( data39                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[39]  )
    );

    idu_rf_preg idu_rf_preg40(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[40]            ),
        .write_data     ( write_data40            ),
        .data           ( data40                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[40]  )
    );

    idu_rf_preg idu_rf_preg41(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[41]            ),
        .write_data     ( write_data41            ),
        .data           ( data41                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[41]  )
    );

    idu_rf_preg idu_rf_preg42(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[42]            ),
        .write_data     ( write_data42            ),
        .data           ( data42                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[42]  )
    );

    idu_rf_preg idu_rf_preg43(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[43]            ),
        .write_data     ( write_data43            ),
        .data           ( data43                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[43]  )
    );

    idu_rf_preg idu_rf_preg44(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[44]            ),
        .write_data     ( write_data44            ),
        .data           ( data44                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[44]  )
    );

    idu_rf_preg idu_rf_preg45(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[45]            ),
        .write_data     ( write_data45            ),
        .data           ( data45                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[45]  )
    );

    idu_rf_preg idu_rf_preg46(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[46]            ),
        .write_data     ( write_data46            ),
        .data           ( data46                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[46]  )
    );

    idu_rf_preg idu_rf_preg47(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[47]            ),
        .write_data     ( write_data47            ),
        .data           ( data47                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[47]  )
    );

    idu_rf_preg idu_rf_preg48(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[48]            ),
        .write_data     ( write_data48            ),
        .data           ( data48                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[48]  )
    );

    idu_rf_preg idu_rf_preg49(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[49]            ),
        .write_data     ( write_data49            ),
        .data           ( data49                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[49]  )
    );

    idu_rf_preg idu_rf_preg50(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[50]            ),
        .write_data     ( write_data50            ),
        .data           ( data50                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[50]  )
    );

    idu_rf_preg idu_rf_preg51(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[51]            ),
        .write_data     ( write_data51            ),
        .data           ( data51                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[51]  )
    );

    idu_rf_preg idu_rf_preg52(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[52]            ),
        .write_data     ( write_data52            ),
        .data           ( data52                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[52]  )
    );

    idu_rf_preg idu_rf_preg53(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[53]            ),
        .write_data     ( write_data53            ),
        .data           ( data53                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[53]  )
    );

    idu_rf_preg idu_rf_preg54(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[54]            ),
        .write_data     ( write_data54            ),
        .data           ( data54                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[54]  )
    );

    idu_rf_preg idu_rf_preg55(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[55]            ),
        .write_data     ( write_data55            ),
        .data           ( data55                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[55]  )
    );

    idu_rf_preg idu_rf_preg56(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[56]            ),
        .write_data     ( write_data56            ),
        .data           ( data56                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[56]  )
    );

    idu_rf_preg idu_rf_preg57(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[57]            ),
        .write_data     ( write_data57            ),
        .data           ( data57                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[57]  )
    );

    idu_rf_preg idu_rf_preg58(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[58]            ),
        .write_data     ( write_data58            ),
        .data           ( data58                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[58]  )
    );

    idu_rf_preg idu_rf_preg59(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[59]            ),
        .write_data     ( write_data59            ),
        .data           ( data59                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[59]  )
    );

    idu_rf_preg idu_rf_preg60(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[60]            ),
        .write_data     ( write_data60            ),
        .data           ( data60                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[60]  )
    );

    idu_rf_preg idu_rf_preg61(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[61]            ),
        .write_data     ( write_data61            ),
        .data           ( data61                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[61]  )
    );

    idu_rf_preg idu_rf_preg62(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[62]            ),
        .write_data     ( write_data62            ),
        .data           ( data62                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[62]  )
    );

    idu_rf_preg idu_rf_preg63(
        .clk            ( clk                    ),
        .rst_clk        ( rst_clk                ),
        .write_en       ( write_en[63]            ),
        .write_data     ( write_data63            ),
        .data           ( data63                  ),
        .wb_vld         ( idu_rtu_pst_wb_vld[63]  )
    );

    assign pipe0_psrc1_decode[0]  = (idu_idu_rf_x_pipe0_psrc1 == 6'd0 );
    assign pipe0_psrc1_decode[1]  = (idu_idu_rf_x_pipe0_psrc1 == 6'd1 );
    assign pipe0_psrc1_decode[2]  = (idu_idu_rf_x_pipe0_psrc1 == 6'd2 );
    assign pipe0_psrc1_decode[3]  = (idu_idu_rf_x_pipe0_psrc1 == 6'd3 );
    assign pipe0_psrc1_decode[4]  = (idu_idu_rf_x_pipe0_psrc1 == 6'd4 );
    assign pipe0_psrc1_decode[5]  = (idu_idu_rf_x_pipe0_psrc1 == 6'd5 );
    assign pipe0_psrc1_decode[6]  = (idu_idu_rf_x_pipe0_psrc1 == 6'd6 );
    assign pipe0_psrc1_decode[7]  = (idu_idu_rf_x_pipe0_psrc1 == 6'd7 );
    assign pipe0_psrc1_decode[8]  = (idu_idu_rf_x_pipe0_psrc1 == 6'd8 );
    assign pipe0_psrc1_decode[9]  = (idu_idu_rf_x_pipe0_psrc1 == 6'd9 );
    assign pipe0_psrc1_decode[10] = (idu_idu_rf_x_pipe0_psrc1 == 6'd10);
    assign pipe0_psrc1_decode[11] = (idu_idu_rf_x_pipe0_psrc1 == 6'd11);
    assign pipe0_psrc1_decode[12] = (idu_idu_rf_x_pipe0_psrc1 == 6'd12);
    assign pipe0_psrc1_decode[13] = (idu_idu_rf_x_pipe0_psrc1 == 6'd13);
    assign pipe0_psrc1_decode[14] = (idu_idu_rf_x_pipe0_psrc1 == 6'd14);
    assign pipe0_psrc1_decode[15] = (idu_idu_rf_x_pipe0_psrc1 == 6'd15);
    assign pipe0_psrc1_decode[16] = (idu_idu_rf_x_pipe0_psrc1 == 6'd16);
    assign pipe0_psrc1_decode[17] = (idu_idu_rf_x_pipe0_psrc1 == 6'd17);
    assign pipe0_psrc1_decode[18] = (idu_idu_rf_x_pipe0_psrc1 == 6'd18);
    assign pipe0_psrc1_decode[19] = (idu_idu_rf_x_pipe0_psrc1 == 6'd19);
    assign pipe0_psrc1_decode[20] = (idu_idu_rf_x_pipe0_psrc1 == 6'd20);
    assign pipe0_psrc1_decode[21] = (idu_idu_rf_x_pipe0_psrc1 == 6'd21);
    assign pipe0_psrc1_decode[22] = (idu_idu_rf_x_pipe0_psrc1 == 6'd22);
    assign pipe0_psrc1_decode[23] = (idu_idu_rf_x_pipe0_psrc1 == 6'd23);
    assign pipe0_psrc1_decode[24] = (idu_idu_rf_x_pipe0_psrc1 == 6'd24);
    assign pipe0_psrc1_decode[25] = (idu_idu_rf_x_pipe0_psrc1 == 6'd25);
    assign pipe0_psrc1_decode[26] = (idu_idu_rf_x_pipe0_psrc1 == 6'd26);
    assign pipe0_psrc1_decode[27] = (idu_idu_rf_x_pipe0_psrc1 == 6'd27);
    assign pipe0_psrc1_decode[28] = (idu_idu_rf_x_pipe0_psrc1 == 6'd28);
    assign pipe0_psrc1_decode[29] = (idu_idu_rf_x_pipe0_psrc1 == 6'd29);
    assign pipe0_psrc1_decode[30] = (idu_idu_rf_x_pipe0_psrc1 == 6'd30);
    assign pipe0_psrc1_decode[31] = (idu_idu_rf_x_pipe0_psrc1 == 6'd31);
    assign pipe0_psrc1_decode[32] = (idu_idu_rf_x_pipe0_psrc1 == 6'd32);
    assign pipe0_psrc1_decode[33] = (idu_idu_rf_x_pipe0_psrc1 == 6'd33);
    assign pipe0_psrc1_decode[34] = (idu_idu_rf_x_pipe0_psrc1 == 6'd34);
    assign pipe0_psrc1_decode[35] = (idu_idu_rf_x_pipe0_psrc1 == 6'd35);
    assign pipe0_psrc1_decode[36] = (idu_idu_rf_x_pipe0_psrc1 == 6'd36);
    assign pipe0_psrc1_decode[37] = (idu_idu_rf_x_pipe0_psrc1 == 6'd37);
    assign pipe0_psrc1_decode[38] = (idu_idu_rf_x_pipe0_psrc1 == 6'd38);
    assign pipe0_psrc1_decode[39] = (idu_idu_rf_x_pipe0_psrc1 == 6'd39);
    assign pipe0_psrc1_decode[40] = (idu_idu_rf_x_pipe0_psrc1 == 6'd40);
    assign pipe0_psrc1_decode[41] = (idu_idu_rf_x_pipe0_psrc1 == 6'd41);
    assign pipe0_psrc1_decode[42] = (idu_idu_rf_x_pipe0_psrc1 == 6'd42);
    assign pipe0_psrc1_decode[43] = (idu_idu_rf_x_pipe0_psrc1 == 6'd43);
    assign pipe0_psrc1_decode[44] = (idu_idu_rf_x_pipe0_psrc1 == 6'd44);
    assign pipe0_psrc1_decode[45] = (idu_idu_rf_x_pipe0_psrc1 == 6'd45);
    assign pipe0_psrc1_decode[46] = (idu_idu_rf_x_pipe0_psrc1 == 6'd46);
    assign pipe0_psrc1_decode[47] = (idu_idu_rf_x_pipe0_psrc1 == 6'd47);
    assign pipe0_psrc1_decode[48] = (idu_idu_rf_x_pipe0_psrc1 == 6'd48);
    assign pipe0_psrc1_decode[49] = (idu_idu_rf_x_pipe0_psrc1 == 6'd49);
    assign pipe0_psrc1_decode[50] = (idu_idu_rf_x_pipe0_psrc1 == 6'd50);
    assign pipe0_psrc1_decode[51] = (idu_idu_rf_x_pipe0_psrc1 == 6'd51);
    assign pipe0_psrc1_decode[52] = (idu_idu_rf_x_pipe0_psrc1 == 6'd52);
    assign pipe0_psrc1_decode[53] = (idu_idu_rf_x_pipe0_psrc1 == 6'd53);
    assign pipe0_psrc1_decode[54] = (idu_idu_rf_x_pipe0_psrc1 == 6'd54);
    assign pipe0_psrc1_decode[55] = (idu_idu_rf_x_pipe0_psrc1 == 6'd55);
    assign pipe0_psrc1_decode[56] = (idu_idu_rf_x_pipe0_psrc1 == 6'd56);
    assign pipe0_psrc1_decode[57] = (idu_idu_rf_x_pipe0_psrc1 == 6'd57);
    assign pipe0_psrc1_decode[58] = (idu_idu_rf_x_pipe0_psrc1 == 6'd58);
    assign pipe0_psrc1_decode[59] = (idu_idu_rf_x_pipe0_psrc1 == 6'd59);
    assign pipe0_psrc1_decode[60] = (idu_idu_rf_x_pipe0_psrc1 == 6'd60);
    assign pipe0_psrc1_decode[61] = (idu_idu_rf_x_pipe0_psrc1 == 6'd61);
    assign pipe0_psrc1_decode[62] = (idu_idu_rf_x_pipe0_psrc1 == 6'd62);
    assign pipe0_psrc1_decode[63] = (idu_idu_rf_x_pipe0_psrc1 == 6'd63);
    assign pipe0_psrc2_decode[0]  = (idu_idu_rf_x_pipe0_psrc2 == 6'd0 );
    assign pipe0_psrc2_decode[1]  = (idu_idu_rf_x_pipe0_psrc2 == 6'd1 );
    assign pipe0_psrc2_decode[2]  = (idu_idu_rf_x_pipe0_psrc2 == 6'd2 );
    assign pipe0_psrc2_decode[3]  = (idu_idu_rf_x_pipe0_psrc2 == 6'd3 );
    assign pipe0_psrc2_decode[4]  = (idu_idu_rf_x_pipe0_psrc2 == 6'd4 );
    assign pipe0_psrc2_decode[5]  = (idu_idu_rf_x_pipe0_psrc2 == 6'd5 );
    assign pipe0_psrc2_decode[6]  = (idu_idu_rf_x_pipe0_psrc2 == 6'd6 );
    assign pipe0_psrc2_decode[7]  = (idu_idu_rf_x_pipe0_psrc2 == 6'd7 );
    assign pipe0_psrc2_decode[8]  = (idu_idu_rf_x_pipe0_psrc2 == 6'd8 );
    assign pipe0_psrc2_decode[9]  = (idu_idu_rf_x_pipe0_psrc2 == 6'd9 );
    assign pipe0_psrc2_decode[10] = (idu_idu_rf_x_pipe0_psrc2 == 6'd10);
    assign pipe0_psrc2_decode[11] = (idu_idu_rf_x_pipe0_psrc2 == 6'd11);
    assign pipe0_psrc2_decode[12] = (idu_idu_rf_x_pipe0_psrc2 == 6'd12);
    assign pipe0_psrc2_decode[13] = (idu_idu_rf_x_pipe0_psrc2 == 6'd13);
    assign pipe0_psrc2_decode[14] = (idu_idu_rf_x_pipe0_psrc2 == 6'd14);
    assign pipe0_psrc2_decode[15] = (idu_idu_rf_x_pipe0_psrc2 == 6'd15);
    assign pipe0_psrc2_decode[16] = (idu_idu_rf_x_pipe0_psrc2 == 6'd16);
    assign pipe0_psrc2_decode[17] = (idu_idu_rf_x_pipe0_psrc2 == 6'd17);
    assign pipe0_psrc2_decode[18] = (idu_idu_rf_x_pipe0_psrc2 == 6'd18);
    assign pipe0_psrc2_decode[19] = (idu_idu_rf_x_pipe0_psrc2 == 6'd19);
    assign pipe0_psrc2_decode[20] = (idu_idu_rf_x_pipe0_psrc2 == 6'd20);
    assign pipe0_psrc2_decode[21] = (idu_idu_rf_x_pipe0_psrc2 == 6'd21);
    assign pipe0_psrc2_decode[22] = (idu_idu_rf_x_pipe0_psrc2 == 6'd22);
    assign pipe0_psrc2_decode[23] = (idu_idu_rf_x_pipe0_psrc2 == 6'd23);
    assign pipe0_psrc2_decode[24] = (idu_idu_rf_x_pipe0_psrc2 == 6'd24);
    assign pipe0_psrc2_decode[25] = (idu_idu_rf_x_pipe0_psrc2 == 6'd25);
    assign pipe0_psrc2_decode[26] = (idu_idu_rf_x_pipe0_psrc2 == 6'd26);
    assign pipe0_psrc2_decode[27] = (idu_idu_rf_x_pipe0_psrc2 == 6'd27);
    assign pipe0_psrc2_decode[28] = (idu_idu_rf_x_pipe0_psrc2 == 6'd28);
    assign pipe0_psrc2_decode[29] = (idu_idu_rf_x_pipe0_psrc2 == 6'd29);
    assign pipe0_psrc2_decode[30] = (idu_idu_rf_x_pipe0_psrc2 == 6'd30);
    assign pipe0_psrc2_decode[31] = (idu_idu_rf_x_pipe0_psrc2 == 6'd31);
    assign pipe0_psrc2_decode[32] = (idu_idu_rf_x_pipe0_psrc2 == 6'd32);
    assign pipe0_psrc2_decode[33] = (idu_idu_rf_x_pipe0_psrc2 == 6'd33);
    assign pipe0_psrc2_decode[34] = (idu_idu_rf_x_pipe0_psrc2 == 6'd34);
    assign pipe0_psrc2_decode[35] = (idu_idu_rf_x_pipe0_psrc2 == 6'd35);
    assign pipe0_psrc2_decode[36] = (idu_idu_rf_x_pipe0_psrc2 == 6'd36);
    assign pipe0_psrc2_decode[37] = (idu_idu_rf_x_pipe0_psrc2 == 6'd37);
    assign pipe0_psrc2_decode[38] = (idu_idu_rf_x_pipe0_psrc2 == 6'd38);
    assign pipe0_psrc2_decode[39] = (idu_idu_rf_x_pipe0_psrc2 == 6'd39);
    assign pipe0_psrc2_decode[40] = (idu_idu_rf_x_pipe0_psrc2 == 6'd40);
    assign pipe0_psrc2_decode[41] = (idu_idu_rf_x_pipe0_psrc2 == 6'd41);
    assign pipe0_psrc2_decode[42] = (idu_idu_rf_x_pipe0_psrc2 == 6'd42);
    assign pipe0_psrc2_decode[43] = (idu_idu_rf_x_pipe0_psrc2 == 6'd43);
    assign pipe0_psrc2_decode[44] = (idu_idu_rf_x_pipe0_psrc2 == 6'd44);
    assign pipe0_psrc2_decode[45] = (idu_idu_rf_x_pipe0_psrc2 == 6'd45);
    assign pipe0_psrc2_decode[46] = (idu_idu_rf_x_pipe0_psrc2 == 6'd46);
    assign pipe0_psrc2_decode[47] = (idu_idu_rf_x_pipe0_psrc2 == 6'd47);
    assign pipe0_psrc2_decode[48] = (idu_idu_rf_x_pipe0_psrc2 == 6'd48);
    assign pipe0_psrc2_decode[49] = (idu_idu_rf_x_pipe0_psrc2 == 6'd49);
    assign pipe0_psrc2_decode[50] = (idu_idu_rf_x_pipe0_psrc2 == 6'd50);
    assign pipe0_psrc2_decode[51] = (idu_idu_rf_x_pipe0_psrc2 == 6'd51);
    assign pipe0_psrc2_decode[52] = (idu_idu_rf_x_pipe0_psrc2 == 6'd52);
    assign pipe0_psrc2_decode[53] = (idu_idu_rf_x_pipe0_psrc2 == 6'd53);
    assign pipe0_psrc2_decode[54] = (idu_idu_rf_x_pipe0_psrc2 == 6'd54);
    assign pipe0_psrc2_decode[55] = (idu_idu_rf_x_pipe0_psrc2 == 6'd55);
    assign pipe0_psrc2_decode[56] = (idu_idu_rf_x_pipe0_psrc2 == 6'd56);
    assign pipe0_psrc2_decode[57] = (idu_idu_rf_x_pipe0_psrc2 == 6'd57);
    assign pipe0_psrc2_decode[58] = (idu_idu_rf_x_pipe0_psrc2 == 6'd58);
    assign pipe0_psrc2_decode[59] = (idu_idu_rf_x_pipe0_psrc2 == 6'd59);
    assign pipe0_psrc2_decode[60] = (idu_idu_rf_x_pipe0_psrc2 == 6'd60);
    assign pipe0_psrc2_decode[61] = (idu_idu_rf_x_pipe0_psrc2 == 6'd61);
    assign pipe0_psrc2_decode[62] = (idu_idu_rf_x_pipe0_psrc2 == 6'd62);
    assign pipe0_psrc2_decode[63] = (idu_idu_rf_x_pipe0_psrc2 == 6'd63);

    assign pipe1_psrc1_decode[0]  = (idu_idu_rf_x_pipe1_psrc1 == 6'd0 );
    assign pipe1_psrc1_decode[1]  = (idu_idu_rf_x_pipe1_psrc1 == 6'd1 );
    assign pipe1_psrc1_decode[2]  = (idu_idu_rf_x_pipe1_psrc1 == 6'd2 );
    assign pipe1_psrc1_decode[3]  = (idu_idu_rf_x_pipe1_psrc1 == 6'd3 );
    assign pipe1_psrc1_decode[4]  = (idu_idu_rf_x_pipe1_psrc1 == 6'd4 );
    assign pipe1_psrc1_decode[5]  = (idu_idu_rf_x_pipe1_psrc1 == 6'd5 );
    assign pipe1_psrc1_decode[6]  = (idu_idu_rf_x_pipe1_psrc1 == 6'd6 );
    assign pipe1_psrc1_decode[7]  = (idu_idu_rf_x_pipe1_psrc1 == 6'd7 );
    assign pipe1_psrc1_decode[8]  = (idu_idu_rf_x_pipe1_psrc1 == 6'd8 );
    assign pipe1_psrc1_decode[9]  = (idu_idu_rf_x_pipe1_psrc1 == 6'd9 );
    assign pipe1_psrc1_decode[10] = (idu_idu_rf_x_pipe1_psrc1 == 6'd10);
    assign pipe1_psrc1_decode[11] = (idu_idu_rf_x_pipe1_psrc1 == 6'd11);
    assign pipe1_psrc1_decode[12] = (idu_idu_rf_x_pipe1_psrc1 == 6'd12);
    assign pipe1_psrc1_decode[13] = (idu_idu_rf_x_pipe1_psrc1 == 6'd13);
    assign pipe1_psrc1_decode[14] = (idu_idu_rf_x_pipe1_psrc1 == 6'd14);
    assign pipe1_psrc1_decode[15] = (idu_idu_rf_x_pipe1_psrc1 == 6'd15);
    assign pipe1_psrc1_decode[16] = (idu_idu_rf_x_pipe1_psrc1 == 6'd16);
    assign pipe1_psrc1_decode[17] = (idu_idu_rf_x_pipe1_psrc1 == 6'd17);
    assign pipe1_psrc1_decode[18] = (idu_idu_rf_x_pipe1_psrc1 == 6'd18);
    assign pipe1_psrc1_decode[19] = (idu_idu_rf_x_pipe1_psrc1 == 6'd19);
    assign pipe1_psrc1_decode[20] = (idu_idu_rf_x_pipe1_psrc1 == 6'd20);
    assign pipe1_psrc1_decode[21] = (idu_idu_rf_x_pipe1_psrc1 == 6'd21);
    assign pipe1_psrc1_decode[22] = (idu_idu_rf_x_pipe1_psrc1 == 6'd22);
    assign pipe1_psrc1_decode[23] = (idu_idu_rf_x_pipe1_psrc1 == 6'd23);
    assign pipe1_psrc1_decode[24] = (idu_idu_rf_x_pipe1_psrc1 == 6'd24);
    assign pipe1_psrc1_decode[25] = (idu_idu_rf_x_pipe1_psrc1 == 6'd25);
    assign pipe1_psrc1_decode[26] = (idu_idu_rf_x_pipe1_psrc1 == 6'd26);
    assign pipe1_psrc1_decode[27] = (idu_idu_rf_x_pipe1_psrc1 == 6'd27);
    assign pipe1_psrc1_decode[28] = (idu_idu_rf_x_pipe1_psrc1 == 6'd28);
    assign pipe1_psrc1_decode[29] = (idu_idu_rf_x_pipe1_psrc1 == 6'd29);
    assign pipe1_psrc1_decode[30] = (idu_idu_rf_x_pipe1_psrc1 == 6'd30);
    assign pipe1_psrc1_decode[31] = (idu_idu_rf_x_pipe1_psrc1 == 6'd31);
    assign pipe1_psrc1_decode[32] = (idu_idu_rf_x_pipe1_psrc1 == 6'd32);
    assign pipe1_psrc1_decode[33] = (idu_idu_rf_x_pipe1_psrc1 == 6'd33);
    assign pipe1_psrc1_decode[34] = (idu_idu_rf_x_pipe1_psrc1 == 6'd34);
    assign pipe1_psrc1_decode[35] = (idu_idu_rf_x_pipe1_psrc1 == 6'd35);
    assign pipe1_psrc1_decode[36] = (idu_idu_rf_x_pipe1_psrc1 == 6'd36);
    assign pipe1_psrc1_decode[37] = (idu_idu_rf_x_pipe1_psrc1 == 6'd37);
    assign pipe1_psrc1_decode[38] = (idu_idu_rf_x_pipe1_psrc1 == 6'd38);
    assign pipe1_psrc1_decode[39] = (idu_idu_rf_x_pipe1_psrc1 == 6'd39);
    assign pipe1_psrc1_decode[40] = (idu_idu_rf_x_pipe1_psrc1 == 6'd40);
    assign pipe1_psrc1_decode[41] = (idu_idu_rf_x_pipe1_psrc1 == 6'd41);
    assign pipe1_psrc1_decode[42] = (idu_idu_rf_x_pipe1_psrc1 == 6'd42);
    assign pipe1_psrc1_decode[43] = (idu_idu_rf_x_pipe1_psrc1 == 6'd43);
    assign pipe1_psrc1_decode[44] = (idu_idu_rf_x_pipe1_psrc1 == 6'd44);
    assign pipe1_psrc1_decode[45] = (idu_idu_rf_x_pipe1_psrc1 == 6'd45);
    assign pipe1_psrc1_decode[46] = (idu_idu_rf_x_pipe1_psrc1 == 6'd46);
    assign pipe1_psrc1_decode[47] = (idu_idu_rf_x_pipe1_psrc1 == 6'd47);
    assign pipe1_psrc1_decode[48] = (idu_idu_rf_x_pipe1_psrc1 == 6'd48);
    assign pipe1_psrc1_decode[49] = (idu_idu_rf_x_pipe1_psrc1 == 6'd49);
    assign pipe1_psrc1_decode[50] = (idu_idu_rf_x_pipe1_psrc1 == 6'd50);
    assign pipe1_psrc1_decode[51] = (idu_idu_rf_x_pipe1_psrc1 == 6'd51);
    assign pipe1_psrc1_decode[52] = (idu_idu_rf_x_pipe1_psrc1 == 6'd52);
    assign pipe1_psrc1_decode[53] = (idu_idu_rf_x_pipe1_psrc1 == 6'd53);
    assign pipe1_psrc1_decode[54] = (idu_idu_rf_x_pipe1_psrc1 == 6'd54);
    assign pipe1_psrc1_decode[55] = (idu_idu_rf_x_pipe1_psrc1 == 6'd55);
    assign pipe1_psrc1_decode[56] = (idu_idu_rf_x_pipe1_psrc1 == 6'd56);
    assign pipe1_psrc1_decode[57] = (idu_idu_rf_x_pipe1_psrc1 == 6'd57);
    assign pipe1_psrc1_decode[58] = (idu_idu_rf_x_pipe1_psrc1 == 6'd58);
    assign pipe1_psrc1_decode[59] = (idu_idu_rf_x_pipe1_psrc1 == 6'd59);
    assign pipe1_psrc1_decode[60] = (idu_idu_rf_x_pipe1_psrc1 == 6'd60);
    assign pipe1_psrc1_decode[61] = (idu_idu_rf_x_pipe1_psrc1 == 6'd61);
    assign pipe1_psrc1_decode[62] = (idu_idu_rf_x_pipe1_psrc1 == 6'd62);
    assign pipe1_psrc1_decode[63] = (idu_idu_rf_x_pipe1_psrc1 == 6'd63);
    assign pipe1_psrc2_decode[0]  = (idu_idu_rf_x_pipe1_psrc2 == 6'd0 );
    assign pipe1_psrc2_decode[1]  = (idu_idu_rf_x_pipe1_psrc2 == 6'd1 );
    assign pipe1_psrc2_decode[2]  = (idu_idu_rf_x_pipe1_psrc2 == 6'd2 );
    assign pipe1_psrc2_decode[3]  = (idu_idu_rf_x_pipe1_psrc2 == 6'd3 );
    assign pipe1_psrc2_decode[4]  = (idu_idu_rf_x_pipe1_psrc2 == 6'd4 );
    assign pipe1_psrc2_decode[5]  = (idu_idu_rf_x_pipe1_psrc2 == 6'd5 );
    assign pipe1_psrc2_decode[6]  = (idu_idu_rf_x_pipe1_psrc2 == 6'd6 );
    assign pipe1_psrc2_decode[7]  = (idu_idu_rf_x_pipe1_psrc2 == 6'd7 );
    assign pipe1_psrc2_decode[8]  = (idu_idu_rf_x_pipe1_psrc2 == 6'd8 );
    assign pipe1_psrc2_decode[9]  = (idu_idu_rf_x_pipe1_psrc2 == 6'd9 );
    assign pipe1_psrc2_decode[10] = (idu_idu_rf_x_pipe1_psrc2 == 6'd10);
    assign pipe1_psrc2_decode[11] = (idu_idu_rf_x_pipe1_psrc2 == 6'd11);
    assign pipe1_psrc2_decode[12] = (idu_idu_rf_x_pipe1_psrc2 == 6'd12);
    assign pipe1_psrc2_decode[13] = (idu_idu_rf_x_pipe1_psrc2 == 6'd13);
    assign pipe1_psrc2_decode[14] = (idu_idu_rf_x_pipe1_psrc2 == 6'd14);
    assign pipe1_psrc2_decode[15] = (idu_idu_rf_x_pipe1_psrc2 == 6'd15);
    assign pipe1_psrc2_decode[16] = (idu_idu_rf_x_pipe1_psrc2 == 6'd16);
    assign pipe1_psrc2_decode[17] = (idu_idu_rf_x_pipe1_psrc2 == 6'd17);
    assign pipe1_psrc2_decode[18] = (idu_idu_rf_x_pipe1_psrc2 == 6'd18);
    assign pipe1_psrc2_decode[19] = (idu_idu_rf_x_pipe1_psrc2 == 6'd19);
    assign pipe1_psrc2_decode[20] = (idu_idu_rf_x_pipe1_psrc2 == 6'd20);
    assign pipe1_psrc2_decode[21] = (idu_idu_rf_x_pipe1_psrc2 == 6'd21);
    assign pipe1_psrc2_decode[22] = (idu_idu_rf_x_pipe1_psrc2 == 6'd22);
    assign pipe1_psrc2_decode[23] = (idu_idu_rf_x_pipe1_psrc2 == 6'd23);
    assign pipe1_psrc2_decode[24] = (idu_idu_rf_x_pipe1_psrc2 == 6'd24);
    assign pipe1_psrc2_decode[25] = (idu_idu_rf_x_pipe1_psrc2 == 6'd25);
    assign pipe1_psrc2_decode[26] = (idu_idu_rf_x_pipe1_psrc2 == 6'd26);
    assign pipe1_psrc2_decode[27] = (idu_idu_rf_x_pipe1_psrc2 == 6'd27);
    assign pipe1_psrc2_decode[28] = (idu_idu_rf_x_pipe1_psrc2 == 6'd28);
    assign pipe1_psrc2_decode[29] = (idu_idu_rf_x_pipe1_psrc2 == 6'd29);
    assign pipe1_psrc2_decode[30] = (idu_idu_rf_x_pipe1_psrc2 == 6'd30);
    assign pipe1_psrc2_decode[31] = (idu_idu_rf_x_pipe1_psrc2 == 6'd31);
    assign pipe1_psrc2_decode[32] = (idu_idu_rf_x_pipe1_psrc2 == 6'd32);
    assign pipe1_psrc2_decode[33] = (idu_idu_rf_x_pipe1_psrc2 == 6'd33);
    assign pipe1_psrc2_decode[34] = (idu_idu_rf_x_pipe1_psrc2 == 6'd34);
    assign pipe1_psrc2_decode[35] = (idu_idu_rf_x_pipe1_psrc2 == 6'd35);
    assign pipe1_psrc2_decode[36] = (idu_idu_rf_x_pipe1_psrc2 == 6'd36);
    assign pipe1_psrc2_decode[37] = (idu_idu_rf_x_pipe1_psrc2 == 6'd37);
    assign pipe1_psrc2_decode[38] = (idu_idu_rf_x_pipe1_psrc2 == 6'd38);
    assign pipe1_psrc2_decode[39] = (idu_idu_rf_x_pipe1_psrc2 == 6'd39);
    assign pipe1_psrc2_decode[40] = (idu_idu_rf_x_pipe1_psrc2 == 6'd40);
    assign pipe1_psrc2_decode[41] = (idu_idu_rf_x_pipe1_psrc2 == 6'd41);
    assign pipe1_psrc2_decode[42] = (idu_idu_rf_x_pipe1_psrc2 == 6'd42);
    assign pipe1_psrc2_decode[43] = (idu_idu_rf_x_pipe1_psrc2 == 6'd43);
    assign pipe1_psrc2_decode[44] = (idu_idu_rf_x_pipe1_psrc2 == 6'd44);
    assign pipe1_psrc2_decode[45] = (idu_idu_rf_x_pipe1_psrc2 == 6'd45);
    assign pipe1_psrc2_decode[46] = (idu_idu_rf_x_pipe1_psrc2 == 6'd46);
    assign pipe1_psrc2_decode[47] = (idu_idu_rf_x_pipe1_psrc2 == 6'd47);
    assign pipe1_psrc2_decode[48] = (idu_idu_rf_x_pipe1_psrc2 == 6'd48);
    assign pipe1_psrc2_decode[49] = (idu_idu_rf_x_pipe1_psrc2 == 6'd49);
    assign pipe1_psrc2_decode[50] = (idu_idu_rf_x_pipe1_psrc2 == 6'd50);
    assign pipe1_psrc2_decode[51] = (idu_idu_rf_x_pipe1_psrc2 == 6'd51);
    assign pipe1_psrc2_decode[52] = (idu_idu_rf_x_pipe1_psrc2 == 6'd52);
    assign pipe1_psrc2_decode[53] = (idu_idu_rf_x_pipe1_psrc2 == 6'd53);
    assign pipe1_psrc2_decode[54] = (idu_idu_rf_x_pipe1_psrc2 == 6'd54);
    assign pipe1_psrc2_decode[55] = (idu_idu_rf_x_pipe1_psrc2 == 6'd55);
    assign pipe1_psrc2_decode[56] = (idu_idu_rf_x_pipe1_psrc2 == 6'd56);
    assign pipe1_psrc2_decode[57] = (idu_idu_rf_x_pipe1_psrc2 == 6'd57);
    assign pipe1_psrc2_decode[58] = (idu_idu_rf_x_pipe1_psrc2 == 6'd58);
    assign pipe1_psrc2_decode[59] = (idu_idu_rf_x_pipe1_psrc2 == 6'd59);
    assign pipe1_psrc2_decode[60] = (idu_idu_rf_x_pipe1_psrc2 == 6'd60);
    assign pipe1_psrc2_decode[61] = (idu_idu_rf_x_pipe1_psrc2 == 6'd61);
    assign pipe1_psrc2_decode[62] = (idu_idu_rf_x_pipe1_psrc2 == 6'd62);
    assign pipe1_psrc2_decode[63] = (idu_idu_rf_x_pipe1_psrc2 == 6'd63);

    assign pipe2_psrc1_decode[0]  = (idu_idu_rf_x_pipe2_psrc1 == 6'd0 );
    assign pipe2_psrc1_decode[1]  = (idu_idu_rf_x_pipe2_psrc1 == 6'd1 );
    assign pipe2_psrc1_decode[2]  = (idu_idu_rf_x_pipe2_psrc1 == 6'd2 );
    assign pipe2_psrc1_decode[3]  = (idu_idu_rf_x_pipe2_psrc1 == 6'd3 );
    assign pipe2_psrc1_decode[4]  = (idu_idu_rf_x_pipe2_psrc1 == 6'd4 );
    assign pipe2_psrc1_decode[5]  = (idu_idu_rf_x_pipe2_psrc1 == 6'd5 );
    assign pipe2_psrc1_decode[6]  = (idu_idu_rf_x_pipe2_psrc1 == 6'd6 );
    assign pipe2_psrc1_decode[7]  = (idu_idu_rf_x_pipe2_psrc1 == 6'd7 );
    assign pipe2_psrc1_decode[8]  = (idu_idu_rf_x_pipe2_psrc1 == 6'd8 );
    assign pipe2_psrc1_decode[9]  = (idu_idu_rf_x_pipe2_psrc1 == 6'd9 );
    assign pipe2_psrc1_decode[10] = (idu_idu_rf_x_pipe2_psrc1 == 6'd10);
    assign pipe2_psrc1_decode[11] = (idu_idu_rf_x_pipe2_psrc1 == 6'd11);
    assign pipe2_psrc1_decode[12] = (idu_idu_rf_x_pipe2_psrc1 == 6'd12);
    assign pipe2_psrc1_decode[13] = (idu_idu_rf_x_pipe2_psrc1 == 6'd13);
    assign pipe2_psrc1_decode[14] = (idu_idu_rf_x_pipe2_psrc1 == 6'd14);
    assign pipe2_psrc1_decode[15] = (idu_idu_rf_x_pipe2_psrc1 == 6'd15);
    assign pipe2_psrc1_decode[16] = (idu_idu_rf_x_pipe2_psrc1 == 6'd16);
    assign pipe2_psrc1_decode[17] = (idu_idu_rf_x_pipe2_psrc1 == 6'd17);
    assign pipe2_psrc1_decode[18] = (idu_idu_rf_x_pipe2_psrc1 == 6'd18);
    assign pipe2_psrc1_decode[19] = (idu_idu_rf_x_pipe2_psrc1 == 6'd19);
    assign pipe2_psrc1_decode[20] = (idu_idu_rf_x_pipe2_psrc1 == 6'd20);
    assign pipe2_psrc1_decode[21] = (idu_idu_rf_x_pipe2_psrc1 == 6'd21);
    assign pipe2_psrc1_decode[22] = (idu_idu_rf_x_pipe2_psrc1 == 6'd22);
    assign pipe2_psrc1_decode[23] = (idu_idu_rf_x_pipe2_psrc1 == 6'd23);
    assign pipe2_psrc1_decode[24] = (idu_idu_rf_x_pipe2_psrc1 == 6'd24);
    assign pipe2_psrc1_decode[25] = (idu_idu_rf_x_pipe2_psrc1 == 6'd25);
    assign pipe2_psrc1_decode[26] = (idu_idu_rf_x_pipe2_psrc1 == 6'd26);
    assign pipe2_psrc1_decode[27] = (idu_idu_rf_x_pipe2_psrc1 == 6'd27);
    assign pipe2_psrc1_decode[28] = (idu_idu_rf_x_pipe2_psrc1 == 6'd28);
    assign pipe2_psrc1_decode[29] = (idu_idu_rf_x_pipe2_psrc1 == 6'd29);
    assign pipe2_psrc1_decode[30] = (idu_idu_rf_x_pipe2_psrc1 == 6'd30);
    assign pipe2_psrc1_decode[31] = (idu_idu_rf_x_pipe2_psrc1 == 6'd31);
    assign pipe2_psrc1_decode[32] = (idu_idu_rf_x_pipe2_psrc1 == 6'd32);
    assign pipe2_psrc1_decode[33] = (idu_idu_rf_x_pipe2_psrc1 == 6'd33);
    assign pipe2_psrc1_decode[34] = (idu_idu_rf_x_pipe2_psrc1 == 6'd34);
    assign pipe2_psrc1_decode[35] = (idu_idu_rf_x_pipe2_psrc1 == 6'd35);
    assign pipe2_psrc1_decode[36] = (idu_idu_rf_x_pipe2_psrc1 == 6'd36);
    assign pipe2_psrc1_decode[37] = (idu_idu_rf_x_pipe2_psrc1 == 6'd37);
    assign pipe2_psrc1_decode[38] = (idu_idu_rf_x_pipe2_psrc1 == 6'd38);
    assign pipe2_psrc1_decode[39] = (idu_idu_rf_x_pipe2_psrc1 == 6'd39);
    assign pipe2_psrc1_decode[40] = (idu_idu_rf_x_pipe2_psrc1 == 6'd40);
    assign pipe2_psrc1_decode[41] = (idu_idu_rf_x_pipe2_psrc1 == 6'd41);
    assign pipe2_psrc1_decode[42] = (idu_idu_rf_x_pipe2_psrc1 == 6'd42);
    assign pipe2_psrc1_decode[43] = (idu_idu_rf_x_pipe2_psrc1 == 6'd43);
    assign pipe2_psrc1_decode[44] = (idu_idu_rf_x_pipe2_psrc1 == 6'd44);
    assign pipe2_psrc1_decode[45] = (idu_idu_rf_x_pipe2_psrc1 == 6'd45);
    assign pipe2_psrc1_decode[46] = (idu_idu_rf_x_pipe2_psrc1 == 6'd46);
    assign pipe2_psrc1_decode[47] = (idu_idu_rf_x_pipe2_psrc1 == 6'd47);
    assign pipe2_psrc1_decode[48] = (idu_idu_rf_x_pipe2_psrc1 == 6'd48);
    assign pipe2_psrc1_decode[49] = (idu_idu_rf_x_pipe2_psrc1 == 6'd49);
    assign pipe2_psrc1_decode[50] = (idu_idu_rf_x_pipe2_psrc1 == 6'd50);
    assign pipe2_psrc1_decode[51] = (idu_idu_rf_x_pipe2_psrc1 == 6'd51);
    assign pipe2_psrc1_decode[52] = (idu_idu_rf_x_pipe2_psrc1 == 6'd52);
    assign pipe2_psrc1_decode[53] = (idu_idu_rf_x_pipe2_psrc1 == 6'd53);
    assign pipe2_psrc1_decode[54] = (idu_idu_rf_x_pipe2_psrc1 == 6'd54);
    assign pipe2_psrc1_decode[55] = (idu_idu_rf_x_pipe2_psrc1 == 6'd55);
    assign pipe2_psrc1_decode[56] = (idu_idu_rf_x_pipe2_psrc1 == 6'd56);
    assign pipe2_psrc1_decode[57] = (idu_idu_rf_x_pipe2_psrc1 == 6'd57);
    assign pipe2_psrc1_decode[58] = (idu_idu_rf_x_pipe2_psrc1 == 6'd58);
    assign pipe2_psrc1_decode[59] = (idu_idu_rf_x_pipe2_psrc1 == 6'd59);
    assign pipe2_psrc1_decode[60] = (idu_idu_rf_x_pipe2_psrc1 == 6'd60);
    assign pipe2_psrc1_decode[61] = (idu_idu_rf_x_pipe2_psrc1 == 6'd61);
    assign pipe2_psrc1_decode[62] = (idu_idu_rf_x_pipe2_psrc1 == 6'd62);
    assign pipe2_psrc1_decode[63] = (idu_idu_rf_x_pipe2_psrc1 == 6'd63);
    assign pipe2_psrc2_decode[0]  = (idu_idu_rf_x_pipe2_psrc2 == 6'd0 );
    assign pipe2_psrc2_decode[1]  = (idu_idu_rf_x_pipe2_psrc2 == 6'd1 );
    assign pipe2_psrc2_decode[2]  = (idu_idu_rf_x_pipe2_psrc2 == 6'd2 );
    assign pipe2_psrc2_decode[3]  = (idu_idu_rf_x_pipe2_psrc2 == 6'd3 );
    assign pipe2_psrc2_decode[4]  = (idu_idu_rf_x_pipe2_psrc2 == 6'd4 );
    assign pipe2_psrc2_decode[5]  = (idu_idu_rf_x_pipe2_psrc2 == 6'd5 );
    assign pipe2_psrc2_decode[6]  = (idu_idu_rf_x_pipe2_psrc2 == 6'd6 );
    assign pipe2_psrc2_decode[7]  = (idu_idu_rf_x_pipe2_psrc2 == 6'd7 );
    assign pipe2_psrc2_decode[8]  = (idu_idu_rf_x_pipe2_psrc2 == 6'd8 );
    assign pipe2_psrc2_decode[9]  = (idu_idu_rf_x_pipe2_psrc2 == 6'd9 );
    assign pipe2_psrc2_decode[10] = (idu_idu_rf_x_pipe2_psrc2 == 6'd10);
    assign pipe2_psrc2_decode[11] = (idu_idu_rf_x_pipe2_psrc2 == 6'd11);
    assign pipe2_psrc2_decode[12] = (idu_idu_rf_x_pipe2_psrc2 == 6'd12);
    assign pipe2_psrc2_decode[13] = (idu_idu_rf_x_pipe2_psrc2 == 6'd13);
    assign pipe2_psrc2_decode[14] = (idu_idu_rf_x_pipe2_psrc2 == 6'd14);
    assign pipe2_psrc2_decode[15] = (idu_idu_rf_x_pipe2_psrc2 == 6'd15);
    assign pipe2_psrc2_decode[16] = (idu_idu_rf_x_pipe2_psrc2 == 6'd16);
    assign pipe2_psrc2_decode[17] = (idu_idu_rf_x_pipe2_psrc2 == 6'd17);
    assign pipe2_psrc2_decode[18] = (idu_idu_rf_x_pipe2_psrc2 == 6'd18);
    assign pipe2_psrc2_decode[19] = (idu_idu_rf_x_pipe2_psrc2 == 6'd19);
    assign pipe2_psrc2_decode[20] = (idu_idu_rf_x_pipe2_psrc2 == 6'd20);
    assign pipe2_psrc2_decode[21] = (idu_idu_rf_x_pipe2_psrc2 == 6'd21);
    assign pipe2_psrc2_decode[22] = (idu_idu_rf_x_pipe2_psrc2 == 6'd22);
    assign pipe2_psrc2_decode[23] = (idu_idu_rf_x_pipe2_psrc2 == 6'd23);
    assign pipe2_psrc2_decode[24] = (idu_idu_rf_x_pipe2_psrc2 == 6'd24);
    assign pipe2_psrc2_decode[25] = (idu_idu_rf_x_pipe2_psrc2 == 6'd25);
    assign pipe2_psrc2_decode[26] = (idu_idu_rf_x_pipe2_psrc2 == 6'd26);
    assign pipe2_psrc2_decode[27] = (idu_idu_rf_x_pipe2_psrc2 == 6'd27);
    assign pipe2_psrc2_decode[28] = (idu_idu_rf_x_pipe2_psrc2 == 6'd28);
    assign pipe2_psrc2_decode[29] = (idu_idu_rf_x_pipe2_psrc2 == 6'd29);
    assign pipe2_psrc2_decode[30] = (idu_idu_rf_x_pipe2_psrc2 == 6'd30);
    assign pipe2_psrc2_decode[31] = (idu_idu_rf_x_pipe2_psrc2 == 6'd31);
    assign pipe2_psrc2_decode[32] = (idu_idu_rf_x_pipe2_psrc2 == 6'd32);
    assign pipe2_psrc2_decode[33] = (idu_idu_rf_x_pipe2_psrc2 == 6'd33);
    assign pipe2_psrc2_decode[34] = (idu_idu_rf_x_pipe2_psrc2 == 6'd34);
    assign pipe2_psrc2_decode[35] = (idu_idu_rf_x_pipe2_psrc2 == 6'd35);
    assign pipe2_psrc2_decode[36] = (idu_idu_rf_x_pipe2_psrc2 == 6'd36);
    assign pipe2_psrc2_decode[37] = (idu_idu_rf_x_pipe2_psrc2 == 6'd37);
    assign pipe2_psrc2_decode[38] = (idu_idu_rf_x_pipe2_psrc2 == 6'd38);
    assign pipe2_psrc2_decode[39] = (idu_idu_rf_x_pipe2_psrc2 == 6'd39);
    assign pipe2_psrc2_decode[40] = (idu_idu_rf_x_pipe2_psrc2 == 6'd40);
    assign pipe2_psrc2_decode[41] = (idu_idu_rf_x_pipe2_psrc2 == 6'd41);
    assign pipe2_psrc2_decode[42] = (idu_idu_rf_x_pipe2_psrc2 == 6'd42);
    assign pipe2_psrc2_decode[43] = (idu_idu_rf_x_pipe2_psrc2 == 6'd43);
    assign pipe2_psrc2_decode[44] = (idu_idu_rf_x_pipe2_psrc2 == 6'd44);
    assign pipe2_psrc2_decode[45] = (idu_idu_rf_x_pipe2_psrc2 == 6'd45);
    assign pipe2_psrc2_decode[46] = (idu_idu_rf_x_pipe2_psrc2 == 6'd46);
    assign pipe2_psrc2_decode[47] = (idu_idu_rf_x_pipe2_psrc2 == 6'd47);
    assign pipe2_psrc2_decode[48] = (idu_idu_rf_x_pipe2_psrc2 == 6'd48);
    assign pipe2_psrc2_decode[49] = (idu_idu_rf_x_pipe2_psrc2 == 6'd49);
    assign pipe2_psrc2_decode[50] = (idu_idu_rf_x_pipe2_psrc2 == 6'd50);
    assign pipe2_psrc2_decode[51] = (idu_idu_rf_x_pipe2_psrc2 == 6'd51);
    assign pipe2_psrc2_decode[52] = (idu_idu_rf_x_pipe2_psrc2 == 6'd52);
    assign pipe2_psrc2_decode[53] = (idu_idu_rf_x_pipe2_psrc2 == 6'd53);
    assign pipe2_psrc2_decode[54] = (idu_idu_rf_x_pipe2_psrc2 == 6'd54);
    assign pipe2_psrc2_decode[55] = (idu_idu_rf_x_pipe2_psrc2 == 6'd55);
    assign pipe2_psrc2_decode[56] = (idu_idu_rf_x_pipe2_psrc2 == 6'd56);
    assign pipe2_psrc2_decode[57] = (idu_idu_rf_x_pipe2_psrc2 == 6'd57);
    assign pipe2_psrc2_decode[58] = (idu_idu_rf_x_pipe2_psrc2 == 6'd58);
    assign pipe2_psrc2_decode[59] = (idu_idu_rf_x_pipe2_psrc2 == 6'd59);
    assign pipe2_psrc2_decode[60] = (idu_idu_rf_x_pipe2_psrc2 == 6'd60);
    assign pipe2_psrc2_decode[61] = (idu_idu_rf_x_pipe2_psrc2 == 6'd61);
    assign pipe2_psrc2_decode[62] = (idu_idu_rf_x_pipe2_psrc2 == 6'd62);
    assign pipe2_psrc2_decode[63] = (idu_idu_rf_x_pipe2_psrc2 == 6'd63);

    assign pipe3_psrc1_decode[0]  = (idu_idu_rf_x_pipe3_psrc1 == 6'd0 );
    assign pipe3_psrc1_decode[1]  = (idu_idu_rf_x_pipe3_psrc1 == 6'd1 );
    assign pipe3_psrc1_decode[2]  = (idu_idu_rf_x_pipe3_psrc1 == 6'd2 );
    assign pipe3_psrc1_decode[3]  = (idu_idu_rf_x_pipe3_psrc1 == 6'd3 );
    assign pipe3_psrc1_decode[4]  = (idu_idu_rf_x_pipe3_psrc1 == 6'd4 );
    assign pipe3_psrc1_decode[5]  = (idu_idu_rf_x_pipe3_psrc1 == 6'd5 );
    assign pipe3_psrc1_decode[6]  = (idu_idu_rf_x_pipe3_psrc1 == 6'd6 );
    assign pipe3_psrc1_decode[7]  = (idu_idu_rf_x_pipe3_psrc1 == 6'd7 );
    assign pipe3_psrc1_decode[8]  = (idu_idu_rf_x_pipe3_psrc1 == 6'd8 );
    assign pipe3_psrc1_decode[9]  = (idu_idu_rf_x_pipe3_psrc1 == 6'd9 );
    assign pipe3_psrc1_decode[10] = (idu_idu_rf_x_pipe3_psrc1 == 6'd10);
    assign pipe3_psrc1_decode[11] = (idu_idu_rf_x_pipe3_psrc1 == 6'd11);
    assign pipe3_psrc1_decode[12] = (idu_idu_rf_x_pipe3_psrc1 == 6'd12);
    assign pipe3_psrc1_decode[13] = (idu_idu_rf_x_pipe3_psrc1 == 6'd13);
    assign pipe3_psrc1_decode[14] = (idu_idu_rf_x_pipe3_psrc1 == 6'd14);
    assign pipe3_psrc1_decode[15] = (idu_idu_rf_x_pipe3_psrc1 == 6'd15);
    assign pipe3_psrc1_decode[16] = (idu_idu_rf_x_pipe3_psrc1 == 6'd16);
    assign pipe3_psrc1_decode[17] = (idu_idu_rf_x_pipe3_psrc1 == 6'd17);
    assign pipe3_psrc1_decode[18] = (idu_idu_rf_x_pipe3_psrc1 == 6'd18);
    assign pipe3_psrc1_decode[19] = (idu_idu_rf_x_pipe3_psrc1 == 6'd19);
    assign pipe3_psrc1_decode[20] = (idu_idu_rf_x_pipe3_psrc1 == 6'd20);
    assign pipe3_psrc1_decode[21] = (idu_idu_rf_x_pipe3_psrc1 == 6'd21);
    assign pipe3_psrc1_decode[22] = (idu_idu_rf_x_pipe3_psrc1 == 6'd22);
    assign pipe3_psrc1_decode[23] = (idu_idu_rf_x_pipe3_psrc1 == 6'd23);
    assign pipe3_psrc1_decode[24] = (idu_idu_rf_x_pipe3_psrc1 == 6'd24);
    assign pipe3_psrc1_decode[25] = (idu_idu_rf_x_pipe3_psrc1 == 6'd25);
    assign pipe3_psrc1_decode[26] = (idu_idu_rf_x_pipe3_psrc1 == 6'd26);
    assign pipe3_psrc1_decode[27] = (idu_idu_rf_x_pipe3_psrc1 == 6'd27);
    assign pipe3_psrc1_decode[28] = (idu_idu_rf_x_pipe3_psrc1 == 6'd28);
    assign pipe3_psrc1_decode[29] = (idu_idu_rf_x_pipe3_psrc1 == 6'd29);
    assign pipe3_psrc1_decode[30] = (idu_idu_rf_x_pipe3_psrc1 == 6'd30);
    assign pipe3_psrc1_decode[31] = (idu_idu_rf_x_pipe3_psrc1 == 6'd31);
    assign pipe3_psrc1_decode[32] = (idu_idu_rf_x_pipe3_psrc1 == 6'd32);
    assign pipe3_psrc1_decode[33] = (idu_idu_rf_x_pipe3_psrc1 == 6'd33);
    assign pipe3_psrc1_decode[34] = (idu_idu_rf_x_pipe3_psrc1 == 6'd34);
    assign pipe3_psrc1_decode[35] = (idu_idu_rf_x_pipe3_psrc1 == 6'd35);
    assign pipe3_psrc1_decode[36] = (idu_idu_rf_x_pipe3_psrc1 == 6'd36);
    assign pipe3_psrc1_decode[37] = (idu_idu_rf_x_pipe3_psrc1 == 6'd37);
    assign pipe3_psrc1_decode[38] = (idu_idu_rf_x_pipe3_psrc1 == 6'd38);
    assign pipe3_psrc1_decode[39] = (idu_idu_rf_x_pipe3_psrc1 == 6'd39);
    assign pipe3_psrc1_decode[40] = (idu_idu_rf_x_pipe3_psrc1 == 6'd40);
    assign pipe3_psrc1_decode[41] = (idu_idu_rf_x_pipe3_psrc1 == 6'd41);
    assign pipe3_psrc1_decode[42] = (idu_idu_rf_x_pipe3_psrc1 == 6'd42);
    assign pipe3_psrc1_decode[43] = (idu_idu_rf_x_pipe3_psrc1 == 6'd43);
    assign pipe3_psrc1_decode[44] = (idu_idu_rf_x_pipe3_psrc1 == 6'd44);
    assign pipe3_psrc1_decode[45] = (idu_idu_rf_x_pipe3_psrc1 == 6'd45);
    assign pipe3_psrc1_decode[46] = (idu_idu_rf_x_pipe3_psrc1 == 6'd46);
    assign pipe3_psrc1_decode[47] = (idu_idu_rf_x_pipe3_psrc1 == 6'd47);
    assign pipe3_psrc1_decode[48] = (idu_idu_rf_x_pipe3_psrc1 == 6'd48);
    assign pipe3_psrc1_decode[49] = (idu_idu_rf_x_pipe3_psrc1 == 6'd49);
    assign pipe3_psrc1_decode[50] = (idu_idu_rf_x_pipe3_psrc1 == 6'd50);
    assign pipe3_psrc1_decode[51] = (idu_idu_rf_x_pipe3_psrc1 == 6'd51);
    assign pipe3_psrc1_decode[52] = (idu_idu_rf_x_pipe3_psrc1 == 6'd52);
    assign pipe3_psrc1_decode[53] = (idu_idu_rf_x_pipe3_psrc1 == 6'd53);
    assign pipe3_psrc1_decode[54] = (idu_idu_rf_x_pipe3_psrc1 == 6'd54);
    assign pipe3_psrc1_decode[55] = (idu_idu_rf_x_pipe3_psrc1 == 6'd55);
    assign pipe3_psrc1_decode[56] = (idu_idu_rf_x_pipe3_psrc1 == 6'd56);
    assign pipe3_psrc1_decode[57] = (idu_idu_rf_x_pipe3_psrc1 == 6'd57);
    assign pipe3_psrc1_decode[58] = (idu_idu_rf_x_pipe3_psrc1 == 6'd58);
    assign pipe3_psrc1_decode[59] = (idu_idu_rf_x_pipe3_psrc1 == 6'd59);
    assign pipe3_psrc1_decode[60] = (idu_idu_rf_x_pipe3_psrc1 == 6'd60);
    assign pipe3_psrc1_decode[61] = (idu_idu_rf_x_pipe3_psrc1 == 6'd61);
    assign pipe3_psrc1_decode[62] = (idu_idu_rf_x_pipe3_psrc1 == 6'd62);
    assign pipe3_psrc1_decode[63] = (idu_idu_rf_x_pipe3_psrc1 == 6'd63);
    assign pipe3_psrc2_decode[0]  = (idu_idu_rf_x_pipe3_psrc2 == 6'd0 );
    assign pipe3_psrc2_decode[1]  = (idu_idu_rf_x_pipe3_psrc2 == 6'd1 );
    assign pipe3_psrc2_decode[2]  = (idu_idu_rf_x_pipe3_psrc2 == 6'd2 );
    assign pipe3_psrc2_decode[3]  = (idu_idu_rf_x_pipe3_psrc2 == 6'd3 );
    assign pipe3_psrc2_decode[4]  = (idu_idu_rf_x_pipe3_psrc2 == 6'd4 );
    assign pipe3_psrc2_decode[5]  = (idu_idu_rf_x_pipe3_psrc2 == 6'd5 );
    assign pipe3_psrc2_decode[6]  = (idu_idu_rf_x_pipe3_psrc2 == 6'd6 );
    assign pipe3_psrc2_decode[7]  = (idu_idu_rf_x_pipe3_psrc2 == 6'd7 );
    assign pipe3_psrc2_decode[8]  = (idu_idu_rf_x_pipe3_psrc2 == 6'd8 );
    assign pipe3_psrc2_decode[9]  = (idu_idu_rf_x_pipe3_psrc2 == 6'd9 );
    assign pipe3_psrc2_decode[10] = (idu_idu_rf_x_pipe3_psrc2 == 6'd10);
    assign pipe3_psrc2_decode[11] = (idu_idu_rf_x_pipe3_psrc2 == 6'd11);
    assign pipe3_psrc2_decode[12] = (idu_idu_rf_x_pipe3_psrc2 == 6'd12);
    assign pipe3_psrc2_decode[13] = (idu_idu_rf_x_pipe3_psrc2 == 6'd13);
    assign pipe3_psrc2_decode[14] = (idu_idu_rf_x_pipe3_psrc2 == 6'd14);
    assign pipe3_psrc2_decode[15] = (idu_idu_rf_x_pipe3_psrc2 == 6'd15);
    assign pipe3_psrc2_decode[16] = (idu_idu_rf_x_pipe3_psrc2 == 6'd16);
    assign pipe3_psrc2_decode[17] = (idu_idu_rf_x_pipe3_psrc2 == 6'd17);
    assign pipe3_psrc2_decode[18] = (idu_idu_rf_x_pipe3_psrc2 == 6'd18);
    assign pipe3_psrc2_decode[19] = (idu_idu_rf_x_pipe3_psrc2 == 6'd19);
    assign pipe3_psrc2_decode[20] = (idu_idu_rf_x_pipe3_psrc2 == 6'd20);
    assign pipe3_psrc2_decode[21] = (idu_idu_rf_x_pipe3_psrc2 == 6'd21);
    assign pipe3_psrc2_decode[22] = (idu_idu_rf_x_pipe3_psrc2 == 6'd22);
    assign pipe3_psrc2_decode[23] = (idu_idu_rf_x_pipe3_psrc2 == 6'd23);
    assign pipe3_psrc2_decode[24] = (idu_idu_rf_x_pipe3_psrc2 == 6'd24);
    assign pipe3_psrc2_decode[25] = (idu_idu_rf_x_pipe3_psrc2 == 6'd25);
    assign pipe3_psrc2_decode[26] = (idu_idu_rf_x_pipe3_psrc2 == 6'd26);
    assign pipe3_psrc2_decode[27] = (idu_idu_rf_x_pipe3_psrc2 == 6'd27);
    assign pipe3_psrc2_decode[28] = (idu_idu_rf_x_pipe3_psrc2 == 6'd28);
    assign pipe3_psrc2_decode[29] = (idu_idu_rf_x_pipe3_psrc2 == 6'd29);
    assign pipe3_psrc2_decode[30] = (idu_idu_rf_x_pipe3_psrc2 == 6'd30);
    assign pipe3_psrc2_decode[31] = (idu_idu_rf_x_pipe3_psrc2 == 6'd31);
    assign pipe3_psrc2_decode[32] = (idu_idu_rf_x_pipe3_psrc2 == 6'd32);
    assign pipe3_psrc2_decode[33] = (idu_idu_rf_x_pipe3_psrc2 == 6'd33);
    assign pipe3_psrc2_decode[34] = (idu_idu_rf_x_pipe3_psrc2 == 6'd34);
    assign pipe3_psrc2_decode[35] = (idu_idu_rf_x_pipe3_psrc2 == 6'd35);
    assign pipe3_psrc2_decode[36] = (idu_idu_rf_x_pipe3_psrc2 == 6'd36);
    assign pipe3_psrc2_decode[37] = (idu_idu_rf_x_pipe3_psrc2 == 6'd37);
    assign pipe3_psrc2_decode[38] = (idu_idu_rf_x_pipe3_psrc2 == 6'd38);
    assign pipe3_psrc2_decode[39] = (idu_idu_rf_x_pipe3_psrc2 == 6'd39);
    assign pipe3_psrc2_decode[40] = (idu_idu_rf_x_pipe3_psrc2 == 6'd40);
    assign pipe3_psrc2_decode[41] = (idu_idu_rf_x_pipe3_psrc2 == 6'd41);
    assign pipe3_psrc2_decode[42] = (idu_idu_rf_x_pipe3_psrc2 == 6'd42);
    assign pipe3_psrc2_decode[43] = (idu_idu_rf_x_pipe3_psrc2 == 6'd43);
    assign pipe3_psrc2_decode[44] = (idu_idu_rf_x_pipe3_psrc2 == 6'd44);
    assign pipe3_psrc2_decode[45] = (idu_idu_rf_x_pipe3_psrc2 == 6'd45);
    assign pipe3_psrc2_decode[46] = (idu_idu_rf_x_pipe3_psrc2 == 6'd46);
    assign pipe3_psrc2_decode[47] = (idu_idu_rf_x_pipe3_psrc2 == 6'd47);
    assign pipe3_psrc2_decode[48] = (idu_idu_rf_x_pipe3_psrc2 == 6'd48);
    assign pipe3_psrc2_decode[49] = (idu_idu_rf_x_pipe3_psrc2 == 6'd49);
    assign pipe3_psrc2_decode[50] = (idu_idu_rf_x_pipe3_psrc2 == 6'd50);
    assign pipe3_psrc2_decode[51] = (idu_idu_rf_x_pipe3_psrc2 == 6'd51);
    assign pipe3_psrc2_decode[52] = (idu_idu_rf_x_pipe3_psrc2 == 6'd52);
    assign pipe3_psrc2_decode[53] = (idu_idu_rf_x_pipe3_psrc2 == 6'd53);
    assign pipe3_psrc2_decode[54] = (idu_idu_rf_x_pipe3_psrc2 == 6'd54);
    assign pipe3_psrc2_decode[55] = (idu_idu_rf_x_pipe3_psrc2 == 6'd55);
    assign pipe3_psrc2_decode[56] = (idu_idu_rf_x_pipe3_psrc2 == 6'd56);
    assign pipe3_psrc2_decode[57] = (idu_idu_rf_x_pipe3_psrc2 == 6'd57);
    assign pipe3_psrc2_decode[58] = (idu_idu_rf_x_pipe3_psrc2 == 6'd58);
    assign pipe3_psrc2_decode[59] = (idu_idu_rf_x_pipe3_psrc2 == 6'd59);
    assign pipe3_psrc2_decode[60] = (idu_idu_rf_x_pipe3_psrc2 == 6'd60);
    assign pipe3_psrc2_decode[61] = (idu_idu_rf_x_pipe3_psrc2 == 6'd61);
    assign pipe3_psrc2_decode[62] = (idu_idu_rf_x_pipe3_psrc2 == 6'd62);
    assign pipe3_psrc2_decode[63] = (idu_idu_rf_x_pipe3_psrc2 == 6'd63);

    assign pipe4_psrc1_decode[0]  = (idu_idu_rf_x_pipe4_psrc1 == 6'd0 );
    assign pipe4_psrc1_decode[1]  = (idu_idu_rf_x_pipe4_psrc1 == 6'd1 );
    assign pipe4_psrc1_decode[2]  = (idu_idu_rf_x_pipe4_psrc1 == 6'd2 );
    assign pipe4_psrc1_decode[3]  = (idu_idu_rf_x_pipe4_psrc1 == 6'd3 );
    assign pipe4_psrc1_decode[4]  = (idu_idu_rf_x_pipe4_psrc1 == 6'd4 );
    assign pipe4_psrc1_decode[5]  = (idu_idu_rf_x_pipe4_psrc1 == 6'd5 );
    assign pipe4_psrc1_decode[6]  = (idu_idu_rf_x_pipe4_psrc1 == 6'd6 );
    assign pipe4_psrc1_decode[7]  = (idu_idu_rf_x_pipe4_psrc1 == 6'd7 );
    assign pipe4_psrc1_decode[8]  = (idu_idu_rf_x_pipe4_psrc1 == 6'd8 );
    assign pipe4_psrc1_decode[9]  = (idu_idu_rf_x_pipe4_psrc1 == 6'd9 );
    assign pipe4_psrc1_decode[10] = (idu_idu_rf_x_pipe4_psrc1 == 6'd10);
    assign pipe4_psrc1_decode[11] = (idu_idu_rf_x_pipe4_psrc1 == 6'd11);
    assign pipe4_psrc1_decode[12] = (idu_idu_rf_x_pipe4_psrc1 == 6'd12);
    assign pipe4_psrc1_decode[13] = (idu_idu_rf_x_pipe4_psrc1 == 6'd13);
    assign pipe4_psrc1_decode[14] = (idu_idu_rf_x_pipe4_psrc1 == 6'd14);
    assign pipe4_psrc1_decode[15] = (idu_idu_rf_x_pipe4_psrc1 == 6'd15);
    assign pipe4_psrc1_decode[16] = (idu_idu_rf_x_pipe4_psrc1 == 6'd16);
    assign pipe4_psrc1_decode[17] = (idu_idu_rf_x_pipe4_psrc1 == 6'd17);
    assign pipe4_psrc1_decode[18] = (idu_idu_rf_x_pipe4_psrc1 == 6'd18);
    assign pipe4_psrc1_decode[19] = (idu_idu_rf_x_pipe4_psrc1 == 6'd19);
    assign pipe4_psrc1_decode[20] = (idu_idu_rf_x_pipe4_psrc1 == 6'd20);
    assign pipe4_psrc1_decode[21] = (idu_idu_rf_x_pipe4_psrc1 == 6'd21);
    assign pipe4_psrc1_decode[22] = (idu_idu_rf_x_pipe4_psrc1 == 6'd22);
    assign pipe4_psrc1_decode[23] = (idu_idu_rf_x_pipe4_psrc1 == 6'd23);
    assign pipe4_psrc1_decode[24] = (idu_idu_rf_x_pipe4_psrc1 == 6'd24);
    assign pipe4_psrc1_decode[25] = (idu_idu_rf_x_pipe4_psrc1 == 6'd25);
    assign pipe4_psrc1_decode[26] = (idu_idu_rf_x_pipe4_psrc1 == 6'd26);
    assign pipe4_psrc1_decode[27] = (idu_idu_rf_x_pipe4_psrc1 == 6'd27);
    assign pipe4_psrc1_decode[28] = (idu_idu_rf_x_pipe4_psrc1 == 6'd28);
    assign pipe4_psrc1_decode[29] = (idu_idu_rf_x_pipe4_psrc1 == 6'd29);
    assign pipe4_psrc1_decode[30] = (idu_idu_rf_x_pipe4_psrc1 == 6'd30);
    assign pipe4_psrc1_decode[31] = (idu_idu_rf_x_pipe4_psrc1 == 6'd31);
    assign pipe4_psrc1_decode[32] = (idu_idu_rf_x_pipe4_psrc1 == 6'd32);
    assign pipe4_psrc1_decode[33] = (idu_idu_rf_x_pipe4_psrc1 == 6'd33);
    assign pipe4_psrc1_decode[34] = (idu_idu_rf_x_pipe4_psrc1 == 6'd34);
    assign pipe4_psrc1_decode[35] = (idu_idu_rf_x_pipe4_psrc1 == 6'd35);
    assign pipe4_psrc1_decode[36] = (idu_idu_rf_x_pipe4_psrc1 == 6'd36);
    assign pipe4_psrc1_decode[37] = (idu_idu_rf_x_pipe4_psrc1 == 6'd37);
    assign pipe4_psrc1_decode[38] = (idu_idu_rf_x_pipe4_psrc1 == 6'd38);
    assign pipe4_psrc1_decode[39] = (idu_idu_rf_x_pipe4_psrc1 == 6'd39);
    assign pipe4_psrc1_decode[40] = (idu_idu_rf_x_pipe4_psrc1 == 6'd40);
    assign pipe4_psrc1_decode[41] = (idu_idu_rf_x_pipe4_psrc1 == 6'd41);
    assign pipe4_psrc1_decode[42] = (idu_idu_rf_x_pipe4_psrc1 == 6'd42);
    assign pipe4_psrc1_decode[43] = (idu_idu_rf_x_pipe4_psrc1 == 6'd43);
    assign pipe4_psrc1_decode[44] = (idu_idu_rf_x_pipe4_psrc1 == 6'd44);
    assign pipe4_psrc1_decode[45] = (idu_idu_rf_x_pipe4_psrc1 == 6'd45);
    assign pipe4_psrc1_decode[46] = (idu_idu_rf_x_pipe4_psrc1 == 6'd46);
    assign pipe4_psrc1_decode[47] = (idu_idu_rf_x_pipe4_psrc1 == 6'd47);
    assign pipe4_psrc1_decode[48] = (idu_idu_rf_x_pipe4_psrc1 == 6'd48);
    assign pipe4_psrc1_decode[49] = (idu_idu_rf_x_pipe4_psrc1 == 6'd49);
    assign pipe4_psrc1_decode[50] = (idu_idu_rf_x_pipe4_psrc1 == 6'd50);
    assign pipe4_psrc1_decode[51] = (idu_idu_rf_x_pipe4_psrc1 == 6'd51);
    assign pipe4_psrc1_decode[52] = (idu_idu_rf_x_pipe4_psrc1 == 6'd52);
    assign pipe4_psrc1_decode[53] = (idu_idu_rf_x_pipe4_psrc1 == 6'd53);
    assign pipe4_psrc1_decode[54] = (idu_idu_rf_x_pipe4_psrc1 == 6'd54);
    assign pipe4_psrc1_decode[55] = (idu_idu_rf_x_pipe4_psrc1 == 6'd55);
    assign pipe4_psrc1_decode[56] = (idu_idu_rf_x_pipe4_psrc1 == 6'd56);
    assign pipe4_psrc1_decode[57] = (idu_idu_rf_x_pipe4_psrc1 == 6'd57);
    assign pipe4_psrc1_decode[58] = (idu_idu_rf_x_pipe4_psrc1 == 6'd58);
    assign pipe4_psrc1_decode[59] = (idu_idu_rf_x_pipe4_psrc1 == 6'd59);
    assign pipe4_psrc1_decode[60] = (idu_idu_rf_x_pipe4_psrc1 == 6'd60);
    assign pipe4_psrc1_decode[61] = (idu_idu_rf_x_pipe4_psrc1 == 6'd61);
    assign pipe4_psrc1_decode[62] = (idu_idu_rf_x_pipe4_psrc1 == 6'd62);
    assign pipe4_psrc1_decode[63] = (idu_idu_rf_x_pipe4_psrc1 == 6'd63);

    // read
    assign idu_idu_rf_x_pipe0_psrc1_value = (idu_idu_rf_x_pipe0_psrc1_vld) ? (
                                                  (data0  & {64{pipe0_psrc1_decode[0]}})
                                                | (data1  & {64{pipe0_psrc1_decode[1]}})
                                                | (data2  & {64{pipe0_psrc1_decode[2]}})
                                                | (data3  & {64{pipe0_psrc1_decode[3]}})
                                                | (data4  & {64{pipe0_psrc1_decode[4]}})
                                                | (data5  & {64{pipe0_psrc1_decode[5]}})
                                                | (data6  & {64{pipe0_psrc1_decode[6]}})
                                                | (data7  & {64{pipe0_psrc1_decode[7]}})
                                                | (data8  & {64{pipe0_psrc1_decode[8]}})
                                                | (data9  & {64{pipe0_psrc1_decode[9]}})
                                                | (data10 & {64{pipe0_psrc1_decode[10]}})
                                                | (data11 & {64{pipe0_psrc1_decode[11]}})
                                                | (data12 & {64{pipe0_psrc1_decode[12]}})
                                                | (data13 & {64{pipe0_psrc1_decode[13]}})
                                                | (data14 & {64{pipe0_psrc1_decode[14]}})
                                                | (data15 & {64{pipe0_psrc1_decode[15]}})
                                                | (data16 & {64{pipe0_psrc1_decode[16]}})
                                                | (data17 & {64{pipe0_psrc1_decode[17]}})
                                                | (data18 & {64{pipe0_psrc1_decode[18]}})
                                                | (data19 & {64{pipe0_psrc1_decode[19]}})
                                                | (data20 & {64{pipe0_psrc1_decode[20]}})
                                                | (data21 & {64{pipe0_psrc1_decode[21]}})
                                                | (data22 & {64{pipe0_psrc1_decode[22]}})
                                                | (data23 & {64{pipe0_psrc1_decode[23]}})
                                                | (data24 & {64{pipe0_psrc1_decode[24]}})
                                                | (data25 & {64{pipe0_psrc1_decode[25]}})
                                                | (data26 & {64{pipe0_psrc1_decode[26]}})
                                                | (data27 & {64{pipe0_psrc1_decode[27]}})
                                                | (data28 & {64{pipe0_psrc1_decode[28]}})
                                                | (data29 & {64{pipe0_psrc1_decode[29]}})
                                                | (data30 & {64{pipe0_psrc1_decode[30]}})
                                                | (data31 & {64{pipe0_psrc1_decode[31]}})
                                                | (data32 & {64{pipe0_psrc1_decode[32]}})
                                                | (data33 & {64{pipe0_psrc1_decode[33]}})
                                                | (data34 & {64{pipe0_psrc1_decode[34]}})
                                                | (data35 & {64{pipe0_psrc1_decode[35]}})
                                                | (data36 & {64{pipe0_psrc1_decode[36]}})
                                                | (data37 & {64{pipe0_psrc1_decode[37]}})
                                                | (data38 & {64{pipe0_psrc1_decode[38]}})
                                                | (data39 & {64{pipe0_psrc1_decode[39]}})
                                                | (data40 & {64{pipe0_psrc1_decode[40]}})
                                                | (data41 & {64{pipe0_psrc1_decode[41]}})
                                                | (data42 & {64{pipe0_psrc1_decode[42]}})
                                                | (data43 & {64{pipe0_psrc1_decode[43]}})
                                                | (data44 & {64{pipe0_psrc1_decode[44]}})
                                                | (data45 & {64{pipe0_psrc1_decode[45]}})
                                                | (data46 & {64{pipe0_psrc1_decode[46]}})
                                                | (data47 & {64{pipe0_psrc1_decode[47]}})
                                                | (data48 & {64{pipe0_psrc1_decode[48]}})
                                                | (data49 & {64{pipe0_psrc1_decode[49]}})
                                                | (data50 & {64{pipe0_psrc1_decode[50]}})
                                                | (data51 & {64{pipe0_psrc1_decode[51]}})
                                                | (data52 & {64{pipe0_psrc1_decode[52]}})
                                                | (data53 & {64{pipe0_psrc1_decode[53]}})
                                                | (data54 & {64{pipe0_psrc1_decode[54]}})
                                                | (data55 & {64{pipe0_psrc1_decode[55]}})
                                                | (data56 & {64{pipe0_psrc1_decode[56]}})
                                                | (data57 & {64{pipe0_psrc1_decode[57]}})
                                                | (data58 & {64{pipe0_psrc1_decode[58]}})
                                                | (data59 & {64{pipe0_psrc1_decode[59]}})
                                                | (data60 & {64{pipe0_psrc1_decode[60]}})
                                                | (data61 & {64{pipe0_psrc1_decode[61]}})
                                                | (data62 & {64{pipe0_psrc1_decode[62]}})
                                                | (data63 & {64{pipe0_psrc1_decode[63]}}))
                                                : 0;
    assign idu_idu_rf_x_pipe0_psrc2_value = (idu_idu_rf_x_pipe0_psrc2_vld) ? (
                                                  (data0  & {64{pipe0_psrc2_decode[0]}})
                                                | (data1  & {64{pipe0_psrc2_decode[1]}})
                                                | (data2  & {64{pipe0_psrc2_decode[2]}})
                                                | (data3  & {64{pipe0_psrc2_decode[3]}})
                                                | (data4  & {64{pipe0_psrc2_decode[4]}})
                                                | (data5  & {64{pipe0_psrc2_decode[5]}})
                                                | (data6  & {64{pipe0_psrc2_decode[6]}})
                                                | (data7  & {64{pipe0_psrc2_decode[7]}})
                                                | (data8  & {64{pipe0_psrc2_decode[8]}})
                                                | (data9  & {64{pipe0_psrc2_decode[9]}})
                                                | (data10 & {64{pipe0_psrc2_decode[10]}})
                                                | (data11 & {64{pipe0_psrc2_decode[11]}})
                                                | (data12 & {64{pipe0_psrc2_decode[12]}})
                                                | (data13 & {64{pipe0_psrc2_decode[13]}})
                                                | (data14 & {64{pipe0_psrc2_decode[14]}})
                                                | (data15 & {64{pipe0_psrc2_decode[15]}})
                                                | (data16 & {64{pipe0_psrc2_decode[16]}})
                                                | (data17 & {64{pipe0_psrc2_decode[17]}})
                                                | (data18 & {64{pipe0_psrc2_decode[18]}})
                                                | (data19 & {64{pipe0_psrc2_decode[19]}})
                                                | (data20 & {64{pipe0_psrc2_decode[20]}})
                                                | (data21 & {64{pipe0_psrc2_decode[21]}})
                                                | (data22 & {64{pipe0_psrc2_decode[22]}})
                                                | (data23 & {64{pipe0_psrc2_decode[23]}})
                                                | (data24 & {64{pipe0_psrc2_decode[24]}})
                                                | (data25 & {64{pipe0_psrc2_decode[25]}})
                                                | (data26 & {64{pipe0_psrc2_decode[26]}})
                                                | (data27 & {64{pipe0_psrc2_decode[27]}})
                                                | (data28 & {64{pipe0_psrc2_decode[28]}})
                                                | (data29 & {64{pipe0_psrc2_decode[29]}})
                                                | (data30 & {64{pipe0_psrc2_decode[30]}})
                                                | (data31 & {64{pipe0_psrc2_decode[31]}})
                                                | (data32 & {64{pipe0_psrc2_decode[32]}})
                                                | (data33 & {64{pipe0_psrc2_decode[33]}})
                                                | (data34 & {64{pipe0_psrc2_decode[34]}})
                                                | (data35 & {64{pipe0_psrc2_decode[35]}})
                                                | (data36 & {64{pipe0_psrc2_decode[36]}})
                                                | (data37 & {64{pipe0_psrc2_decode[37]}})
                                                | (data38 & {64{pipe0_psrc2_decode[38]}})
                                                | (data39 & {64{pipe0_psrc2_decode[39]}})
                                                | (data40 & {64{pipe0_psrc2_decode[40]}})
                                                | (data41 & {64{pipe0_psrc2_decode[41]}})
                                                | (data42 & {64{pipe0_psrc2_decode[42]}})
                                                | (data43 & {64{pipe0_psrc2_decode[43]}})
                                                | (data44 & {64{pipe0_psrc2_decode[44]}})
                                                | (data45 & {64{pipe0_psrc2_decode[45]}})
                                                | (data46 & {64{pipe0_psrc2_decode[46]}})
                                                | (data47 & {64{pipe0_psrc2_decode[47]}})
                                                | (data48 & {64{pipe0_psrc2_decode[48]}})
                                                | (data49 & {64{pipe0_psrc2_decode[49]}})
                                                | (data50 & {64{pipe0_psrc2_decode[50]}})
                                                | (data51 & {64{pipe0_psrc2_decode[51]}})
                                                | (data52 & {64{pipe0_psrc2_decode[52]}})
                                                | (data53 & {64{pipe0_psrc2_decode[53]}})
                                                | (data54 & {64{pipe0_psrc2_decode[54]}})
                                                | (data55 & {64{pipe0_psrc2_decode[55]}})
                                                | (data56 & {64{pipe0_psrc2_decode[56]}})
                                                | (data57 & {64{pipe0_psrc2_decode[57]}})
                                                | (data58 & {64{pipe0_psrc2_decode[58]}})
                                                | (data59 & {64{pipe0_psrc2_decode[59]}})
                                                | (data60 & {64{pipe0_psrc2_decode[60]}})
                                                | (data61 & {64{pipe0_psrc2_decode[61]}})
                                                | (data62 & {64{pipe0_psrc2_decode[62]}})
                                                | (data63 & {64{pipe0_psrc2_decode[63]}}))
                                                : 0;

    assign idu_idu_rf_x_pipe1_psrc1_value = (idu_idu_rf_x_pipe1_psrc1_vld) ? (
                                                  (data0  & {64{pipe1_psrc1_decode[0]}})
                                                | (data1  & {64{pipe1_psrc1_decode[1]}})
                                                | (data2  & {64{pipe1_psrc1_decode[2]}})
                                                | (data3  & {64{pipe1_psrc1_decode[3]}})
                                                | (data4  & {64{pipe1_psrc1_decode[4]}})
                                                | (data5  & {64{pipe1_psrc1_decode[5]}})
                                                | (data6  & {64{pipe1_psrc1_decode[6]}})
                                                | (data7  & {64{pipe1_psrc1_decode[7]}})
                                                | (data8  & {64{pipe1_psrc1_decode[8]}})
                                                | (data9  & {64{pipe1_psrc1_decode[9]}})
                                                | (data10 & {64{pipe1_psrc1_decode[10]}})
                                                | (data11 & {64{pipe1_psrc1_decode[11]}})
                                                | (data12 & {64{pipe1_psrc1_decode[12]}})
                                                | (data13 & {64{pipe1_psrc1_decode[13]}})
                                                | (data14 & {64{pipe1_psrc1_decode[14]}})
                                                | (data15 & {64{pipe1_psrc1_decode[15]}})
                                                | (data16 & {64{pipe1_psrc1_decode[16]}})
                                                | (data17 & {64{pipe1_psrc1_decode[17]}})
                                                | (data18 & {64{pipe1_psrc1_decode[18]}})
                                                | (data19 & {64{pipe1_psrc1_decode[19]}})
                                                | (data20 & {64{pipe1_psrc1_decode[20]}})
                                                | (data21 & {64{pipe1_psrc1_decode[21]}})
                                                | (data22 & {64{pipe1_psrc1_decode[22]}})
                                                | (data23 & {64{pipe1_psrc1_decode[23]}})
                                                | (data24 & {64{pipe1_psrc1_decode[24]}})
                                                | (data25 & {64{pipe1_psrc1_decode[25]}})
                                                | (data26 & {64{pipe1_psrc1_decode[26]}})
                                                | (data27 & {64{pipe1_psrc1_decode[27]}})
                                                | (data28 & {64{pipe1_psrc1_decode[28]}})
                                                | (data29 & {64{pipe1_psrc1_decode[29]}})
                                                | (data30 & {64{pipe1_psrc1_decode[30]}})
                                                | (data31 & {64{pipe1_psrc1_decode[31]}})
                                                | (data32 & {64{pipe1_psrc1_decode[32]}})
                                                | (data33 & {64{pipe1_psrc1_decode[33]}})
                                                | (data34 & {64{pipe1_psrc1_decode[34]}})
                                                | (data35 & {64{pipe1_psrc1_decode[35]}})
                                                | (data36 & {64{pipe1_psrc1_decode[36]}})
                                                | (data37 & {64{pipe1_psrc1_decode[37]}})
                                                | (data38 & {64{pipe1_psrc1_decode[38]}})
                                                | (data39 & {64{pipe1_psrc1_decode[39]}})
                                                | (data40 & {64{pipe1_psrc1_decode[40]}})
                                                | (data41 & {64{pipe1_psrc1_decode[41]}})
                                                | (data42 & {64{pipe1_psrc1_decode[42]}})
                                                | (data43 & {64{pipe1_psrc1_decode[43]}})
                                                | (data44 & {64{pipe1_psrc1_decode[44]}})
                                                | (data45 & {64{pipe1_psrc1_decode[45]}})
                                                | (data46 & {64{pipe1_psrc1_decode[46]}})
                                                | (data47 & {64{pipe1_psrc1_decode[47]}})
                                                | (data48 & {64{pipe1_psrc1_decode[48]}})
                                                | (data49 & {64{pipe1_psrc1_decode[49]}})
                                                | (data50 & {64{pipe1_psrc1_decode[50]}})
                                                | (data51 & {64{pipe1_psrc1_decode[51]}})
                                                | (data52 & {64{pipe1_psrc1_decode[52]}})
                                                | (data53 & {64{pipe1_psrc1_decode[53]}})
                                                | (data54 & {64{pipe1_psrc1_decode[54]}})
                                                | (data55 & {64{pipe1_psrc1_decode[55]}})
                                                | (data56 & {64{pipe1_psrc1_decode[56]}})
                                                | (data57 & {64{pipe1_psrc1_decode[57]}})
                                                | (data58 & {64{pipe1_psrc1_decode[58]}})
                                                | (data59 & {64{pipe1_psrc1_decode[59]}})
                                                | (data60 & {64{pipe1_psrc1_decode[60]}})
                                                | (data61 & {64{pipe1_psrc1_decode[61]}})
                                                | (data62 & {64{pipe1_psrc1_decode[62]}})
                                                | (data63 & {64{pipe1_psrc1_decode[63]}}))
                                                : 0;
    assign idu_idu_rf_x_pipe1_psrc2_value = (idu_idu_rf_x_pipe1_psrc2_vld) ? (
                                                  (data0  & {64{pipe1_psrc2_decode[0]}})
                                                | (data1  & {64{pipe1_psrc2_decode[1]}})
                                                | (data2  & {64{pipe1_psrc2_decode[2]}})
                                                | (data3  & {64{pipe1_psrc2_decode[3]}})
                                                | (data4  & {64{pipe1_psrc2_decode[4]}})
                                                | (data5  & {64{pipe1_psrc2_decode[5]}})
                                                | (data6  & {64{pipe1_psrc2_decode[6]}})
                                                | (data7  & {64{pipe1_psrc2_decode[7]}})
                                                | (data8  & {64{pipe1_psrc2_decode[8]}})
                                                | (data9  & {64{pipe1_psrc2_decode[9]}})
                                                | (data10 & {64{pipe1_psrc2_decode[10]}})
                                                | (data11 & {64{pipe1_psrc2_decode[11]}})
                                                | (data12 & {64{pipe1_psrc2_decode[12]}})
                                                | (data13 & {64{pipe1_psrc2_decode[13]}})
                                                | (data14 & {64{pipe1_psrc2_decode[14]}})
                                                | (data15 & {64{pipe1_psrc2_decode[15]}})
                                                | (data16 & {64{pipe1_psrc2_decode[16]}})
                                                | (data17 & {64{pipe1_psrc2_decode[17]}})
                                                | (data18 & {64{pipe1_psrc2_decode[18]}})
                                                | (data19 & {64{pipe1_psrc2_decode[19]}})
                                                | (data20 & {64{pipe1_psrc2_decode[20]}})
                                                | (data21 & {64{pipe1_psrc2_decode[21]}})
                                                | (data22 & {64{pipe1_psrc2_decode[22]}})
                                                | (data23 & {64{pipe1_psrc2_decode[23]}})
                                                | (data24 & {64{pipe1_psrc2_decode[24]}})
                                                | (data25 & {64{pipe1_psrc2_decode[25]}})
                                                | (data26 & {64{pipe1_psrc2_decode[26]}})
                                                | (data27 & {64{pipe1_psrc2_decode[27]}})
                                                | (data28 & {64{pipe1_psrc2_decode[28]}})
                                                | (data29 & {64{pipe1_psrc2_decode[29]}})
                                                | (data30 & {64{pipe1_psrc2_decode[30]}})
                                                | (data31 & {64{pipe1_psrc2_decode[31]}})
                                                | (data32 & {64{pipe1_psrc2_decode[32]}})
                                                | (data33 & {64{pipe1_psrc2_decode[33]}})
                                                | (data34 & {64{pipe1_psrc2_decode[34]}})
                                                | (data35 & {64{pipe1_psrc2_decode[35]}})
                                                | (data36 & {64{pipe1_psrc2_decode[36]}})
                                                | (data37 & {64{pipe1_psrc2_decode[37]}})
                                                | (data38 & {64{pipe1_psrc2_decode[38]}})
                                                | (data39 & {64{pipe1_psrc2_decode[39]}})
                                                | (data40 & {64{pipe1_psrc2_decode[40]}})
                                                | (data41 & {64{pipe1_psrc2_decode[41]}})
                                                | (data42 & {64{pipe1_psrc2_decode[42]}})
                                                | (data43 & {64{pipe1_psrc2_decode[43]}})
                                                | (data44 & {64{pipe1_psrc2_decode[44]}})
                                                | (data45 & {64{pipe1_psrc2_decode[45]}})
                                                | (data46 & {64{pipe1_psrc2_decode[46]}})
                                                | (data47 & {64{pipe1_psrc2_decode[47]}})
                                                | (data48 & {64{pipe1_psrc2_decode[48]}})
                                                | (data49 & {64{pipe1_psrc2_decode[49]}})
                                                | (data50 & {64{pipe1_psrc2_decode[50]}})
                                                | (data51 & {64{pipe1_psrc2_decode[51]}})
                                                | (data52 & {64{pipe1_psrc2_decode[52]}})
                                                | (data53 & {64{pipe1_psrc2_decode[53]}})
                                                | (data54 & {64{pipe1_psrc2_decode[54]}})
                                                | (data55 & {64{pipe1_psrc2_decode[55]}})
                                                | (data56 & {64{pipe1_psrc2_decode[56]}})
                                                | (data57 & {64{pipe1_psrc2_decode[57]}})
                                                | (data58 & {64{pipe1_psrc2_decode[58]}})
                                                | (data59 & {64{pipe1_psrc2_decode[59]}})
                                                | (data60 & {64{pipe1_psrc2_decode[60]}})
                                                | (data61 & {64{pipe1_psrc2_decode[61]}})
                                                | (data62 & {64{pipe1_psrc2_decode[62]}})
                                                | (data63 & {64{pipe1_psrc2_decode[63]}}))
                                                : 0;

    assign idu_idu_rf_x_pipe2_psrc1_value = (idu_idu_rf_x_pipe2_psrc1_vld) ? (
                                                  (data0  & {64{pipe2_psrc1_decode[0]}})
                                                | (data1  & {64{pipe2_psrc1_decode[1]}})
                                                | (data2  & {64{pipe2_psrc1_decode[2]}})
                                                | (data3  & {64{pipe2_psrc1_decode[3]}})
                                                | (data4  & {64{pipe2_psrc1_decode[4]}})
                                                | (data5  & {64{pipe2_psrc1_decode[5]}})
                                                | (data6  & {64{pipe2_psrc1_decode[6]}})
                                                | (data7  & {64{pipe2_psrc1_decode[7]}})
                                                | (data8  & {64{pipe2_psrc1_decode[8]}})
                                                | (data9  & {64{pipe2_psrc1_decode[9]}})
                                                | (data10 & {64{pipe2_psrc1_decode[10]}})
                                                | (data11 & {64{pipe2_psrc1_decode[11]}})
                                                | (data12 & {64{pipe2_psrc1_decode[12]}})
                                                | (data13 & {64{pipe2_psrc1_decode[13]}})
                                                | (data14 & {64{pipe2_psrc1_decode[14]}})
                                                | (data15 & {64{pipe2_psrc1_decode[15]}})
                                                | (data16 & {64{pipe2_psrc1_decode[16]}})
                                                | (data17 & {64{pipe2_psrc1_decode[17]}})
                                                | (data18 & {64{pipe2_psrc1_decode[18]}})
                                                | (data19 & {64{pipe2_psrc1_decode[19]}})
                                                | (data20 & {64{pipe2_psrc1_decode[20]}})
                                                | (data21 & {64{pipe2_psrc1_decode[21]}})
                                                | (data22 & {64{pipe2_psrc1_decode[22]}})
                                                | (data23 & {64{pipe2_psrc1_decode[23]}})
                                                | (data24 & {64{pipe2_psrc1_decode[24]}})
                                                | (data25 & {64{pipe2_psrc1_decode[25]}})
                                                | (data26 & {64{pipe2_psrc1_decode[26]}})
                                                | (data27 & {64{pipe2_psrc1_decode[27]}})
                                                | (data28 & {64{pipe2_psrc1_decode[28]}})
                                                | (data29 & {64{pipe2_psrc1_decode[29]}})
                                                | (data30 & {64{pipe2_psrc1_decode[30]}})
                                                | (data31 & {64{pipe2_psrc1_decode[31]}})
                                                | (data32 & {64{pipe2_psrc1_decode[32]}})
                                                | (data33 & {64{pipe2_psrc1_decode[33]}})
                                                | (data34 & {64{pipe2_psrc1_decode[34]}})
                                                | (data35 & {64{pipe2_psrc1_decode[35]}})
                                                | (data36 & {64{pipe2_psrc1_decode[36]}})
                                                | (data37 & {64{pipe2_psrc1_decode[37]}})
                                                | (data38 & {64{pipe2_psrc1_decode[38]}})
                                                | (data39 & {64{pipe2_psrc1_decode[39]}})
                                                | (data40 & {64{pipe2_psrc1_decode[40]}})
                                                | (data41 & {64{pipe2_psrc1_decode[41]}})
                                                | (data42 & {64{pipe2_psrc1_decode[42]}})
                                                | (data43 & {64{pipe2_psrc1_decode[43]}})
                                                | (data44 & {64{pipe2_psrc1_decode[44]}})
                                                | (data45 & {64{pipe2_psrc1_decode[45]}})
                                                | (data46 & {64{pipe2_psrc1_decode[46]}})
                                                | (data47 & {64{pipe2_psrc1_decode[47]}})
                                                | (data48 & {64{pipe2_psrc1_decode[48]}})
                                                | (data49 & {64{pipe2_psrc1_decode[49]}})
                                                | (data50 & {64{pipe2_psrc1_decode[50]}})
                                                | (data51 & {64{pipe2_psrc1_decode[51]}})
                                                | (data52 & {64{pipe2_psrc1_decode[52]}})
                                                | (data53 & {64{pipe2_psrc1_decode[53]}})
                                                | (data54 & {64{pipe2_psrc1_decode[54]}})
                                                | (data55 & {64{pipe2_psrc1_decode[55]}})
                                                | (data56 & {64{pipe2_psrc1_decode[56]}})
                                                | (data57 & {64{pipe2_psrc1_decode[57]}})
                                                | (data58 & {64{pipe2_psrc1_decode[58]}})
                                                | (data59 & {64{pipe2_psrc1_decode[59]}})
                                                | (data60 & {64{pipe2_psrc1_decode[60]}})
                                                | (data61 & {64{pipe2_psrc1_decode[61]}})
                                                | (data62 & {64{pipe2_psrc1_decode[62]}})
                                                | (data63 & {64{pipe2_psrc1_decode[63]}}))
                                                : 0;
    assign idu_idu_rf_x_pipe2_psrc2_value = (idu_idu_rf_x_pipe2_psrc2_vld) ? (
                                                  (data0  & {64{pipe2_psrc2_decode[0]}})
                                                | (data1  & {64{pipe2_psrc2_decode[1]}})
                                                | (data2  & {64{pipe2_psrc2_decode[2]}})
                                                | (data3  & {64{pipe2_psrc2_decode[3]}})
                                                | (data4  & {64{pipe2_psrc2_decode[4]}})
                                                | (data5  & {64{pipe2_psrc2_decode[5]}})
                                                | (data6  & {64{pipe2_psrc2_decode[6]}})
                                                | (data7  & {64{pipe2_psrc2_decode[7]}})
                                                | (data8  & {64{pipe2_psrc2_decode[8]}})
                                                | (data9  & {64{pipe2_psrc2_decode[9]}})
                                                | (data10 & {64{pipe2_psrc2_decode[10]}})
                                                | (data11 & {64{pipe2_psrc2_decode[11]}})
                                                | (data12 & {64{pipe2_psrc2_decode[12]}})
                                                | (data13 & {64{pipe2_psrc2_decode[13]}})
                                                | (data14 & {64{pipe2_psrc2_decode[14]}})
                                                | (data15 & {64{pipe2_psrc2_decode[15]}})
                                                | (data16 & {64{pipe2_psrc2_decode[16]}})
                                                | (data17 & {64{pipe2_psrc2_decode[17]}})
                                                | (data18 & {64{pipe2_psrc2_decode[18]}})
                                                | (data19 & {64{pipe2_psrc2_decode[19]}})
                                                | (data20 & {64{pipe2_psrc2_decode[20]}})
                                                | (data21 & {64{pipe2_psrc2_decode[21]}})
                                                | (data22 & {64{pipe2_psrc2_decode[22]}})
                                                | (data23 & {64{pipe2_psrc2_decode[23]}})
                                                | (data24 & {64{pipe2_psrc2_decode[24]}})
                                                | (data25 & {64{pipe2_psrc2_decode[25]}})
                                                | (data26 & {64{pipe2_psrc2_decode[26]}})
                                                | (data27 & {64{pipe2_psrc2_decode[27]}})
                                                | (data28 & {64{pipe2_psrc2_decode[28]}})
                                                | (data29 & {64{pipe2_psrc2_decode[29]}})
                                                | (data30 & {64{pipe2_psrc2_decode[30]}})
                                                | (data31 & {64{pipe2_psrc2_decode[31]}})
                                                | (data32 & {64{pipe2_psrc2_decode[32]}})
                                                | (data33 & {64{pipe2_psrc2_decode[33]}})
                                                | (data34 & {64{pipe2_psrc2_decode[34]}})
                                                | (data35 & {64{pipe2_psrc2_decode[35]}})
                                                | (data36 & {64{pipe2_psrc2_decode[36]}})
                                                | (data37 & {64{pipe2_psrc2_decode[37]}})
                                                | (data38 & {64{pipe2_psrc2_decode[38]}})
                                                | (data39 & {64{pipe2_psrc2_decode[39]}})
                                                | (data40 & {64{pipe2_psrc2_decode[40]}})
                                                | (data41 & {64{pipe2_psrc2_decode[41]}})
                                                | (data42 & {64{pipe2_psrc2_decode[42]}})
                                                | (data43 & {64{pipe2_psrc2_decode[43]}})
                                                | (data44 & {64{pipe2_psrc2_decode[44]}})
                                                | (data45 & {64{pipe2_psrc2_decode[45]}})
                                                | (data46 & {64{pipe2_psrc2_decode[46]}})
                                                | (data47 & {64{pipe2_psrc2_decode[47]}})
                                                | (data48 & {64{pipe2_psrc2_decode[48]}})
                                                | (data49 & {64{pipe2_psrc2_decode[49]}})
                                                | (data50 & {64{pipe2_psrc2_decode[50]}})
                                                | (data51 & {64{pipe2_psrc2_decode[51]}})
                                                | (data52 & {64{pipe2_psrc2_decode[52]}})
                                                | (data53 & {64{pipe2_psrc2_decode[53]}})
                                                | (data54 & {64{pipe2_psrc2_decode[54]}})
                                                | (data55 & {64{pipe2_psrc2_decode[55]}})
                                                | (data56 & {64{pipe2_psrc2_decode[56]}})
                                                | (data57 & {64{pipe2_psrc2_decode[57]}})
                                                | (data58 & {64{pipe2_psrc2_decode[58]}})
                                                | (data59 & {64{pipe2_psrc2_decode[59]}})
                                                | (data60 & {64{pipe2_psrc2_decode[60]}})
                                                | (data61 & {64{pipe2_psrc2_decode[61]}})
                                                | (data62 & {64{pipe2_psrc2_decode[62]}})
                                                | (data63 & {64{pipe2_psrc2_decode[63]}}))
                                                : 0;

    assign idu_idu_rf_x_pipe3_psrc1_value = (idu_idu_rf_x_pipe3_psrc1_vld) ? (
                                                  (data0  & {64{pipe3_psrc1_decode[0]}})
                                                | (data1  & {64{pipe3_psrc1_decode[1]}})
                                                | (data2  & {64{pipe3_psrc1_decode[2]}})
                                                | (data3  & {64{pipe3_psrc1_decode[3]}})
                                                | (data4  & {64{pipe3_psrc1_decode[4]}})
                                                | (data5  & {64{pipe3_psrc1_decode[5]}})
                                                | (data6  & {64{pipe3_psrc1_decode[6]}})
                                                | (data7  & {64{pipe3_psrc1_decode[7]}})
                                                | (data8  & {64{pipe3_psrc1_decode[8]}})
                                                | (data9  & {64{pipe3_psrc1_decode[9]}})
                                                | (data10 & {64{pipe3_psrc1_decode[10]}})
                                                | (data11 & {64{pipe3_psrc1_decode[11]}})
                                                | (data12 & {64{pipe3_psrc1_decode[12]}})
                                                | (data13 & {64{pipe3_psrc1_decode[13]}})
                                                | (data14 & {64{pipe3_psrc1_decode[14]}})
                                                | (data15 & {64{pipe3_psrc1_decode[15]}})
                                                | (data16 & {64{pipe3_psrc1_decode[16]}})
                                                | (data17 & {64{pipe3_psrc1_decode[17]}})
                                                | (data18 & {64{pipe3_psrc1_decode[18]}})
                                                | (data19 & {64{pipe3_psrc1_decode[19]}})
                                                | (data20 & {64{pipe3_psrc1_decode[20]}})
                                                | (data21 & {64{pipe3_psrc1_decode[21]}})
                                                | (data22 & {64{pipe3_psrc1_decode[22]}})
                                                | (data23 & {64{pipe3_psrc1_decode[23]}})
                                                | (data24 & {64{pipe3_psrc1_decode[24]}})
                                                | (data25 & {64{pipe3_psrc1_decode[25]}})
                                                | (data26 & {64{pipe3_psrc1_decode[26]}})
                                                | (data27 & {64{pipe3_psrc1_decode[27]}})
                                                | (data28 & {64{pipe3_psrc1_decode[28]}})
                                                | (data29 & {64{pipe3_psrc1_decode[29]}})
                                                | (data30 & {64{pipe3_psrc1_decode[30]}})
                                                | (data31 & {64{pipe3_psrc1_decode[31]}})
                                                | (data32 & {64{pipe3_psrc1_decode[32]}})
                                                | (data33 & {64{pipe3_psrc1_decode[33]}})
                                                | (data34 & {64{pipe3_psrc1_decode[34]}})
                                                | (data35 & {64{pipe3_psrc1_decode[35]}})
                                                | (data36 & {64{pipe3_psrc1_decode[36]}})
                                                | (data37 & {64{pipe3_psrc1_decode[37]}})
                                                | (data38 & {64{pipe3_psrc1_decode[38]}})
                                                | (data39 & {64{pipe3_psrc1_decode[39]}})
                                                | (data40 & {64{pipe3_psrc1_decode[40]}})
                                                | (data41 & {64{pipe3_psrc1_decode[41]}})
                                                | (data42 & {64{pipe3_psrc1_decode[42]}})
                                                | (data43 & {64{pipe3_psrc1_decode[43]}})
                                                | (data44 & {64{pipe3_psrc1_decode[44]}})
                                                | (data45 & {64{pipe3_psrc1_decode[45]}})
                                                | (data46 & {64{pipe3_psrc1_decode[46]}})
                                                | (data47 & {64{pipe3_psrc1_decode[47]}})
                                                | (data48 & {64{pipe3_psrc1_decode[48]}})
                                                | (data49 & {64{pipe3_psrc1_decode[49]}})
                                                | (data50 & {64{pipe3_psrc1_decode[50]}})
                                                | (data51 & {64{pipe3_psrc1_decode[51]}})
                                                | (data52 & {64{pipe3_psrc1_decode[52]}})
                                                | (data53 & {64{pipe3_psrc1_decode[53]}})
                                                | (data54 & {64{pipe3_psrc1_decode[54]}})
                                                | (data55 & {64{pipe3_psrc1_decode[55]}})
                                                | (data56 & {64{pipe3_psrc1_decode[56]}})
                                                | (data57 & {64{pipe3_psrc1_decode[57]}})
                                                | (data58 & {64{pipe3_psrc1_decode[58]}})
                                                | (data59 & {64{pipe3_psrc1_decode[59]}})
                                                | (data60 & {64{pipe3_psrc1_decode[60]}})
                                                | (data61 & {64{pipe3_psrc1_decode[61]}})
                                                | (data62 & {64{pipe3_psrc1_decode[62]}})
                                                | (data63 & {64{pipe3_psrc1_decode[63]}}))
                                                : 0;
    assign idu_idu_rf_x_pipe3_psrc2_value = (idu_idu_rf_x_pipe3_psrc2_vld) ? (
                                                  (data0  & {64{pipe3_psrc2_decode[0]}})
                                                | (data1  & {64{pipe3_psrc2_decode[1]}})
                                                | (data2  & {64{pipe3_psrc2_decode[2]}})
                                                | (data3  & {64{pipe3_psrc2_decode[3]}})
                                                | (data4  & {64{pipe3_psrc2_decode[4]}})
                                                | (data5  & {64{pipe3_psrc2_decode[5]}})
                                                | (data6  & {64{pipe3_psrc2_decode[6]}})
                                                | (data7  & {64{pipe3_psrc2_decode[7]}})
                                                | (data8  & {64{pipe3_psrc2_decode[8]}})
                                                | (data9  & {64{pipe3_psrc2_decode[9]}})
                                                | (data10 & {64{pipe3_psrc2_decode[10]}})
                                                | (data11 & {64{pipe3_psrc2_decode[11]}})
                                                | (data12 & {64{pipe3_psrc2_decode[12]}})
                                                | (data13 & {64{pipe3_psrc2_decode[13]}})
                                                | (data14 & {64{pipe3_psrc2_decode[14]}})
                                                | (data15 & {64{pipe3_psrc2_decode[15]}})
                                                | (data16 & {64{pipe3_psrc2_decode[16]}})
                                                | (data17 & {64{pipe3_psrc2_decode[17]}})
                                                | (data18 & {64{pipe3_psrc2_decode[18]}})
                                                | (data19 & {64{pipe3_psrc2_decode[19]}})
                                                | (data20 & {64{pipe3_psrc2_decode[20]}})
                                                | (data21 & {64{pipe3_psrc2_decode[21]}})
                                                | (data22 & {64{pipe3_psrc2_decode[22]}})
                                                | (data23 & {64{pipe3_psrc2_decode[23]}})
                                                | (data24 & {64{pipe3_psrc2_decode[24]}})
                                                | (data25 & {64{pipe3_psrc2_decode[25]}})
                                                | (data26 & {64{pipe3_psrc2_decode[26]}})
                                                | (data27 & {64{pipe3_psrc2_decode[27]}})
                                                | (data28 & {64{pipe3_psrc2_decode[28]}})
                                                | (data29 & {64{pipe3_psrc2_decode[29]}})
                                                | (data30 & {64{pipe3_psrc2_decode[30]}})
                                                | (data31 & {64{pipe3_psrc2_decode[31]}})
                                                | (data32 & {64{pipe3_psrc2_decode[32]}})
                                                | (data33 & {64{pipe3_psrc2_decode[33]}})
                                                | (data34 & {64{pipe3_psrc2_decode[34]}})
                                                | (data35 & {64{pipe3_psrc2_decode[35]}})
                                                | (data36 & {64{pipe3_psrc2_decode[36]}})
                                                | (data37 & {64{pipe3_psrc2_decode[37]}})
                                                | (data38 & {64{pipe3_psrc2_decode[38]}})
                                                | (data39 & {64{pipe3_psrc2_decode[39]}})
                                                | (data40 & {64{pipe3_psrc2_decode[40]}})
                                                | (data41 & {64{pipe3_psrc2_decode[41]}})
                                                | (data42 & {64{pipe3_psrc2_decode[42]}})
                                                | (data43 & {64{pipe3_psrc2_decode[43]}})
                                                | (data44 & {64{pipe3_psrc2_decode[44]}})
                                                | (data45 & {64{pipe3_psrc2_decode[45]}})
                                                | (data46 & {64{pipe3_psrc2_decode[46]}})
                                                | (data47 & {64{pipe3_psrc2_decode[47]}})
                                                | (data48 & {64{pipe3_psrc2_decode[48]}})
                                                | (data49 & {64{pipe3_psrc2_decode[49]}})
                                                | (data50 & {64{pipe3_psrc2_decode[50]}})
                                                | (data51 & {64{pipe3_psrc2_decode[51]}})
                                                | (data52 & {64{pipe3_psrc2_decode[52]}})
                                                | (data53 & {64{pipe3_psrc2_decode[53]}})
                                                | (data54 & {64{pipe3_psrc2_decode[54]}})
                                                | (data55 & {64{pipe3_psrc2_decode[55]}})
                                                | (data56 & {64{pipe3_psrc2_decode[56]}})
                                                | (data57 & {64{pipe3_psrc2_decode[57]}})
                                                | (data58 & {64{pipe3_psrc2_decode[58]}})
                                                | (data59 & {64{pipe3_psrc2_decode[59]}})
                                                | (data60 & {64{pipe3_psrc2_decode[60]}})
                                                | (data61 & {64{pipe3_psrc2_decode[61]}})
                                                | (data62 & {64{pipe3_psrc2_decode[62]}})
                                                | (data63 & {64{pipe3_psrc2_decode[63]}}))
                                                : 0;

    assign idu_idu_rf_x_pipe4_psrc1_value = (idu_idu_rf_x_pipe4_psrc1_vld) ? (
                                                  (data0  & {64{pipe4_psrc1_decode[0]}})
                                                | (data1  & {64{pipe4_psrc1_decode[1]}})
                                                | (data2  & {64{pipe4_psrc1_decode[2]}})
                                                | (data3  & {64{pipe4_psrc1_decode[3]}})
                                                | (data4  & {64{pipe4_psrc1_decode[4]}})
                                                | (data5  & {64{pipe4_psrc1_decode[5]}})
                                                | (data6  & {64{pipe4_psrc1_decode[6]}})
                                                | (data7  & {64{pipe4_psrc1_decode[7]}})
                                                | (data8  & {64{pipe4_psrc1_decode[8]}})
                                                | (data9  & {64{pipe4_psrc1_decode[9]}})
                                                | (data10 & {64{pipe4_psrc1_decode[10]}})
                                                | (data11 & {64{pipe4_psrc1_decode[11]}})
                                                | (data12 & {64{pipe4_psrc1_decode[12]}})
                                                | (data13 & {64{pipe4_psrc1_decode[13]}})
                                                | (data14 & {64{pipe4_psrc1_decode[14]}})
                                                | (data15 & {64{pipe4_psrc1_decode[15]}})
                                                | (data16 & {64{pipe4_psrc1_decode[16]}})
                                                | (data17 & {64{pipe4_psrc1_decode[17]}})
                                                | (data18 & {64{pipe4_psrc1_decode[18]}})
                                                | (data19 & {64{pipe4_psrc1_decode[19]}})
                                                | (data20 & {64{pipe4_psrc1_decode[20]}})
                                                | (data21 & {64{pipe4_psrc1_decode[21]}})
                                                | (data22 & {64{pipe4_psrc1_decode[22]}})
                                                | (data23 & {64{pipe4_psrc1_decode[23]}})
                                                | (data24 & {64{pipe4_psrc1_decode[24]}})
                                                | (data25 & {64{pipe4_psrc1_decode[25]}})
                                                | (data26 & {64{pipe4_psrc1_decode[26]}})
                                                | (data27 & {64{pipe4_psrc1_decode[27]}})
                                                | (data28 & {64{pipe4_psrc1_decode[28]}})
                                                | (data29 & {64{pipe4_psrc1_decode[29]}})
                                                | (data30 & {64{pipe4_psrc1_decode[30]}})
                                                | (data31 & {64{pipe4_psrc1_decode[31]}})
                                                | (data32 & {64{pipe4_psrc1_decode[32]}})
                                                | (data33 & {64{pipe4_psrc1_decode[33]}})
                                                | (data34 & {64{pipe4_psrc1_decode[34]}})
                                                | (data35 & {64{pipe4_psrc1_decode[35]}})
                                                | (data36 & {64{pipe4_psrc1_decode[36]}})
                                                | (data37 & {64{pipe4_psrc1_decode[37]}})
                                                | (data38 & {64{pipe4_psrc1_decode[38]}})
                                                | (data39 & {64{pipe4_psrc1_decode[39]}})
                                                | (data40 & {64{pipe4_psrc1_decode[40]}})
                                                | (data41 & {64{pipe4_psrc1_decode[41]}})
                                                | (data42 & {64{pipe4_psrc1_decode[42]}})
                                                | (data43 & {64{pipe4_psrc1_decode[43]}})
                                                | (data44 & {64{pipe4_psrc1_decode[44]}})
                                                | (data45 & {64{pipe4_psrc1_decode[45]}})
                                                | (data46 & {64{pipe4_psrc1_decode[46]}})
                                                | (data47 & {64{pipe4_psrc1_decode[47]}})
                                                | (data48 & {64{pipe4_psrc1_decode[48]}})
                                                | (data49 & {64{pipe4_psrc1_decode[49]}})
                                                | (data50 & {64{pipe4_psrc1_decode[50]}})
                                                | (data51 & {64{pipe4_psrc1_decode[51]}})
                                                | (data52 & {64{pipe4_psrc1_decode[52]}})
                                                | (data53 & {64{pipe4_psrc1_decode[53]}})
                                                | (data54 & {64{pipe4_psrc1_decode[54]}})
                                                | (data55 & {64{pipe4_psrc1_decode[55]}})
                                                | (data56 & {64{pipe4_psrc1_decode[56]}})
                                                | (data57 & {64{pipe4_psrc1_decode[57]}})
                                                | (data58 & {64{pipe4_psrc1_decode[58]}})
                                                | (data59 & {64{pipe4_psrc1_decode[59]}})
                                                | (data60 & {64{pipe4_psrc1_decode[60]}})
                                                | (data61 & {64{pipe4_psrc1_decode[61]}})
                                                | (data62 & {64{pipe4_psrc1_decode[62]}})
                                                | (data63 & {64{pipe4_psrc1_decode[63]}}))
                                                : 0;

    // write
    assign alu_wb_en[0]  = (exu_idu_rf_alu_wb_preg == 6'd0 ) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[1]  = (exu_idu_rf_alu_wb_preg == 6'd1 ) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[2]  = (exu_idu_rf_alu_wb_preg == 6'd2 ) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[3]  = (exu_idu_rf_alu_wb_preg == 6'd3 ) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[4]  = (exu_idu_rf_alu_wb_preg == 6'd4 ) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[5]  = (exu_idu_rf_alu_wb_preg == 6'd5 ) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[6]  = (exu_idu_rf_alu_wb_preg == 6'd6 ) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[7]  = (exu_idu_rf_alu_wb_preg == 6'd7 ) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[8]  = (exu_idu_rf_alu_wb_preg == 6'd8 ) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[9]  = (exu_idu_rf_alu_wb_preg == 6'd9 ) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[10] = (exu_idu_rf_alu_wb_preg == 6'd10) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[11] = (exu_idu_rf_alu_wb_preg == 6'd11) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[12] = (exu_idu_rf_alu_wb_preg == 6'd12) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[13] = (exu_idu_rf_alu_wb_preg == 6'd13) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[14] = (exu_idu_rf_alu_wb_preg == 6'd14) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[15] = (exu_idu_rf_alu_wb_preg == 6'd15) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[16] = (exu_idu_rf_alu_wb_preg == 6'd16) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[17] = (exu_idu_rf_alu_wb_preg == 6'd17) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[18] = (exu_idu_rf_alu_wb_preg == 6'd18) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[19] = (exu_idu_rf_alu_wb_preg == 6'd19) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[20] = (exu_idu_rf_alu_wb_preg == 6'd20) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[21] = (exu_idu_rf_alu_wb_preg == 6'd21) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[22] = (exu_idu_rf_alu_wb_preg == 6'd22) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[23] = (exu_idu_rf_alu_wb_preg == 6'd23) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[24] = (exu_idu_rf_alu_wb_preg == 6'd24) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[25] = (exu_idu_rf_alu_wb_preg == 6'd25) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[26] = (exu_idu_rf_alu_wb_preg == 6'd26) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[27] = (exu_idu_rf_alu_wb_preg == 6'd27) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[28] = (exu_idu_rf_alu_wb_preg == 6'd28) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[29] = (exu_idu_rf_alu_wb_preg == 6'd29) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[30] = (exu_idu_rf_alu_wb_preg == 6'd30) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[31] = (exu_idu_rf_alu_wb_preg == 6'd31) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[32] = (exu_idu_rf_alu_wb_preg == 6'd32) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[33] = (exu_idu_rf_alu_wb_preg == 6'd33) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[34] = (exu_idu_rf_alu_wb_preg == 6'd34) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[35] = (exu_idu_rf_alu_wb_preg == 6'd35) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[36] = (exu_idu_rf_alu_wb_preg == 6'd36) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[37] = (exu_idu_rf_alu_wb_preg == 6'd37) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[38] = (exu_idu_rf_alu_wb_preg == 6'd38) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[39] = (exu_idu_rf_alu_wb_preg == 6'd39) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[40] = (exu_idu_rf_alu_wb_preg == 6'd40) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[41] = (exu_idu_rf_alu_wb_preg == 6'd41) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[42] = (exu_idu_rf_alu_wb_preg == 6'd42) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[43] = (exu_idu_rf_alu_wb_preg == 6'd43) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[44] = (exu_idu_rf_alu_wb_preg == 6'd44) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[45] = (exu_idu_rf_alu_wb_preg == 6'd45) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[46] = (exu_idu_rf_alu_wb_preg == 6'd46) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[47] = (exu_idu_rf_alu_wb_preg == 6'd47) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[48] = (exu_idu_rf_alu_wb_preg == 6'd48) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[49] = (exu_idu_rf_alu_wb_preg == 6'd49) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[50] = (exu_idu_rf_alu_wb_preg == 6'd50) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[51] = (exu_idu_rf_alu_wb_preg == 6'd51) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[52] = (exu_idu_rf_alu_wb_preg == 6'd52) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[53] = (exu_idu_rf_alu_wb_preg == 6'd53) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[54] = (exu_idu_rf_alu_wb_preg == 6'd54) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[55] = (exu_idu_rf_alu_wb_preg == 6'd55) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[56] = (exu_idu_rf_alu_wb_preg == 6'd56) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[57] = (exu_idu_rf_alu_wb_preg == 6'd57) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[58] = (exu_idu_rf_alu_wb_preg == 6'd58) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[59] = (exu_idu_rf_alu_wb_preg == 6'd59) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[60] = (exu_idu_rf_alu_wb_preg == 6'd60) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[61] = (exu_idu_rf_alu_wb_preg == 6'd61) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[62] = (exu_idu_rf_alu_wb_preg == 6'd62) & exu_idu_rf_alu_wb_vld;
    assign alu_wb_en[63] = (exu_idu_rf_alu_wb_preg == 6'd63) & exu_idu_rf_alu_wb_vld;

    assign mxu_wb_en[0]  = (exu_idu_rf_mxu_wb_preg == 6'd0 ) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[1]  = (exu_idu_rf_mxu_wb_preg == 6'd1 ) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[2]  = (exu_idu_rf_mxu_wb_preg == 6'd2 ) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[3]  = (exu_idu_rf_mxu_wb_preg == 6'd3 ) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[4]  = (exu_idu_rf_mxu_wb_preg == 6'd4 ) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[5]  = (exu_idu_rf_mxu_wb_preg == 6'd5 ) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[6]  = (exu_idu_rf_mxu_wb_preg == 6'd6 ) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[7]  = (exu_idu_rf_mxu_wb_preg == 6'd7 ) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[8]  = (exu_idu_rf_mxu_wb_preg == 6'd8 ) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[9]  = (exu_idu_rf_mxu_wb_preg == 6'd9 ) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[10] = (exu_idu_rf_mxu_wb_preg == 6'd10) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[11] = (exu_idu_rf_mxu_wb_preg == 6'd11) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[12] = (exu_idu_rf_mxu_wb_preg == 6'd12) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[13] = (exu_idu_rf_mxu_wb_preg == 6'd13) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[14] = (exu_idu_rf_mxu_wb_preg == 6'd14) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[15] = (exu_idu_rf_mxu_wb_preg == 6'd15) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[16] = (exu_idu_rf_mxu_wb_preg == 6'd16) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[17] = (exu_idu_rf_mxu_wb_preg == 6'd17) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[18] = (exu_idu_rf_mxu_wb_preg == 6'd18) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[19] = (exu_idu_rf_mxu_wb_preg == 6'd19) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[20] = (exu_idu_rf_mxu_wb_preg == 6'd20) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[21] = (exu_idu_rf_mxu_wb_preg == 6'd21) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[22] = (exu_idu_rf_mxu_wb_preg == 6'd22) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[23] = (exu_idu_rf_mxu_wb_preg == 6'd23) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[24] = (exu_idu_rf_mxu_wb_preg == 6'd24) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[25] = (exu_idu_rf_mxu_wb_preg == 6'd25) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[26] = (exu_idu_rf_mxu_wb_preg == 6'd26) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[27] = (exu_idu_rf_mxu_wb_preg == 6'd27) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[28] = (exu_idu_rf_mxu_wb_preg == 6'd28) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[29] = (exu_idu_rf_mxu_wb_preg == 6'd29) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[30] = (exu_idu_rf_mxu_wb_preg == 6'd30) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[31] = (exu_idu_rf_mxu_wb_preg == 6'd31) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[32] = (exu_idu_rf_mxu_wb_preg == 6'd32) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[33] = (exu_idu_rf_mxu_wb_preg == 6'd33) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[34] = (exu_idu_rf_mxu_wb_preg == 6'd34) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[35] = (exu_idu_rf_mxu_wb_preg == 6'd35) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[36] = (exu_idu_rf_mxu_wb_preg == 6'd36) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[37] = (exu_idu_rf_mxu_wb_preg == 6'd37) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[38] = (exu_idu_rf_mxu_wb_preg == 6'd38) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[39] = (exu_idu_rf_mxu_wb_preg == 6'd39) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[40] = (exu_idu_rf_mxu_wb_preg == 6'd40) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[41] = (exu_idu_rf_mxu_wb_preg == 6'd41) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[42] = (exu_idu_rf_mxu_wb_preg == 6'd42) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[43] = (exu_idu_rf_mxu_wb_preg == 6'd43) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[44] = (exu_idu_rf_mxu_wb_preg == 6'd44) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[45] = (exu_idu_rf_mxu_wb_preg == 6'd45) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[46] = (exu_idu_rf_mxu_wb_preg == 6'd46) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[47] = (exu_idu_rf_mxu_wb_preg == 6'd47) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[48] = (exu_idu_rf_mxu_wb_preg == 6'd48) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[49] = (exu_idu_rf_mxu_wb_preg == 6'd49) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[50] = (exu_idu_rf_mxu_wb_preg == 6'd50) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[51] = (exu_idu_rf_mxu_wb_preg == 6'd51) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[52] = (exu_idu_rf_mxu_wb_preg == 6'd52) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[53] = (exu_idu_rf_mxu_wb_preg == 6'd53) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[54] = (exu_idu_rf_mxu_wb_preg == 6'd54) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[55] = (exu_idu_rf_mxu_wb_preg == 6'd55) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[56] = (exu_idu_rf_mxu_wb_preg == 6'd56) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[57] = (exu_idu_rf_mxu_wb_preg == 6'd57) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[58] = (exu_idu_rf_mxu_wb_preg == 6'd58) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[59] = (exu_idu_rf_mxu_wb_preg == 6'd59) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[60] = (exu_idu_rf_mxu_wb_preg == 6'd60) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[61] = (exu_idu_rf_mxu_wb_preg == 6'd61) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[62] = (exu_idu_rf_mxu_wb_preg == 6'd62) & exu_idu_rf_mxu_wb_vld;
    assign mxu_wb_en[63] = (exu_idu_rf_mxu_wb_preg == 6'd63) & exu_idu_rf_mxu_wb_vld;

    assign div_wb_en[0]  = (exu_idu_rf_div_wb_preg == 6'd0 ) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[1]  = (exu_idu_rf_div_wb_preg == 6'd1 ) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[2]  = (exu_idu_rf_div_wb_preg == 6'd2 ) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[3]  = (exu_idu_rf_div_wb_preg == 6'd3 ) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[4]  = (exu_idu_rf_div_wb_preg == 6'd4 ) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[5]  = (exu_idu_rf_div_wb_preg == 6'd5 ) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[6]  = (exu_idu_rf_div_wb_preg == 6'd6 ) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[7]  = (exu_idu_rf_div_wb_preg == 6'd7 ) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[8]  = (exu_idu_rf_div_wb_preg == 6'd8 ) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[9]  = (exu_idu_rf_div_wb_preg == 6'd9 ) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[10] = (exu_idu_rf_div_wb_preg == 6'd10) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[11] = (exu_idu_rf_div_wb_preg == 6'd11) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[12] = (exu_idu_rf_div_wb_preg == 6'd12) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[13] = (exu_idu_rf_div_wb_preg == 6'd13) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[14] = (exu_idu_rf_div_wb_preg == 6'd14) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[15] = (exu_idu_rf_div_wb_preg == 6'd15) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[16] = (exu_idu_rf_div_wb_preg == 6'd16) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[17] = (exu_idu_rf_div_wb_preg == 6'd17) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[18] = (exu_idu_rf_div_wb_preg == 6'd18) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[19] = (exu_idu_rf_div_wb_preg == 6'd19) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[20] = (exu_idu_rf_div_wb_preg == 6'd20) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[21] = (exu_idu_rf_div_wb_preg == 6'd21) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[22] = (exu_idu_rf_div_wb_preg == 6'd22) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[23] = (exu_idu_rf_div_wb_preg == 6'd23) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[24] = (exu_idu_rf_div_wb_preg == 6'd24) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[25] = (exu_idu_rf_div_wb_preg == 6'd25) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[26] = (exu_idu_rf_div_wb_preg == 6'd26) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[27] = (exu_idu_rf_div_wb_preg == 6'd27) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[28] = (exu_idu_rf_div_wb_preg == 6'd28) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[29] = (exu_idu_rf_div_wb_preg == 6'd29) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[30] = (exu_idu_rf_div_wb_preg == 6'd30) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[31] = (exu_idu_rf_div_wb_preg == 6'd31) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[32] = (exu_idu_rf_div_wb_preg == 6'd32) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[33] = (exu_idu_rf_div_wb_preg == 6'd33) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[34] = (exu_idu_rf_div_wb_preg == 6'd34) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[35] = (exu_idu_rf_div_wb_preg == 6'd35) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[36] = (exu_idu_rf_div_wb_preg == 6'd36) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[37] = (exu_idu_rf_div_wb_preg == 6'd37) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[38] = (exu_idu_rf_div_wb_preg == 6'd38) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[39] = (exu_idu_rf_div_wb_preg == 6'd39) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[40] = (exu_idu_rf_div_wb_preg == 6'd40) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[41] = (exu_idu_rf_div_wb_preg == 6'd41) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[42] = (exu_idu_rf_div_wb_preg == 6'd42) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[43] = (exu_idu_rf_div_wb_preg == 6'd43) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[44] = (exu_idu_rf_div_wb_preg == 6'd44) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[45] = (exu_idu_rf_div_wb_preg == 6'd45) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[46] = (exu_idu_rf_div_wb_preg == 6'd46) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[47] = (exu_idu_rf_div_wb_preg == 6'd47) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[48] = (exu_idu_rf_div_wb_preg == 6'd48) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[49] = (exu_idu_rf_div_wb_preg == 6'd49) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[50] = (exu_idu_rf_div_wb_preg == 6'd50) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[51] = (exu_idu_rf_div_wb_preg == 6'd51) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[52] = (exu_idu_rf_div_wb_preg == 6'd52) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[53] = (exu_idu_rf_div_wb_preg == 6'd53) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[54] = (exu_idu_rf_div_wb_preg == 6'd54) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[55] = (exu_idu_rf_div_wb_preg == 6'd55) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[56] = (exu_idu_rf_div_wb_preg == 6'd56) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[57] = (exu_idu_rf_div_wb_preg == 6'd57) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[58] = (exu_idu_rf_div_wb_preg == 6'd58) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[59] = (exu_idu_rf_div_wb_preg == 6'd59) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[60] = (exu_idu_rf_div_wb_preg == 6'd60) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[61] = (exu_idu_rf_div_wb_preg == 6'd61) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[62] = (exu_idu_rf_div_wb_preg == 6'd62) & exu_idu_rf_div_wb_vld;
    assign div_wb_en[63] = (exu_idu_rf_div_wb_preg == 6'd63) & exu_idu_rf_div_wb_vld;

    assign bju_wb_en[0]  = (exu_idu_rf_bju_wb_preg == 6'd0 ) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[1]  = (exu_idu_rf_bju_wb_preg == 6'd1 ) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[2]  = (exu_idu_rf_bju_wb_preg == 6'd2 ) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[3]  = (exu_idu_rf_bju_wb_preg == 6'd3 ) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[4]  = (exu_idu_rf_bju_wb_preg == 6'd4 ) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[5]  = (exu_idu_rf_bju_wb_preg == 6'd5 ) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[6]  = (exu_idu_rf_bju_wb_preg == 6'd6 ) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[7]  = (exu_idu_rf_bju_wb_preg == 6'd7 ) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[8]  = (exu_idu_rf_bju_wb_preg == 6'd8 ) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[9]  = (exu_idu_rf_bju_wb_preg == 6'd9 ) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[10] = (exu_idu_rf_bju_wb_preg == 6'd10) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[11] = (exu_idu_rf_bju_wb_preg == 6'd11) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[12] = (exu_idu_rf_bju_wb_preg == 6'd12) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[13] = (exu_idu_rf_bju_wb_preg == 6'd13) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[14] = (exu_idu_rf_bju_wb_preg == 6'd14) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[15] = (exu_idu_rf_bju_wb_preg == 6'd15) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[16] = (exu_idu_rf_bju_wb_preg == 6'd16) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[17] = (exu_idu_rf_bju_wb_preg == 6'd17) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[18] = (exu_idu_rf_bju_wb_preg == 6'd18) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[19] = (exu_idu_rf_bju_wb_preg == 6'd19) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[20] = (exu_idu_rf_bju_wb_preg == 6'd20) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[21] = (exu_idu_rf_bju_wb_preg == 6'd21) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[22] = (exu_idu_rf_bju_wb_preg == 6'd22) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[23] = (exu_idu_rf_bju_wb_preg == 6'd23) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[24] = (exu_idu_rf_bju_wb_preg == 6'd24) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[25] = (exu_idu_rf_bju_wb_preg == 6'd25) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[26] = (exu_idu_rf_bju_wb_preg == 6'd26) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[27] = (exu_idu_rf_bju_wb_preg == 6'd27) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[28] = (exu_idu_rf_bju_wb_preg == 6'd28) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[29] = (exu_idu_rf_bju_wb_preg == 6'd29) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[30] = (exu_idu_rf_bju_wb_preg == 6'd30) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[31] = (exu_idu_rf_bju_wb_preg == 6'd31) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[32] = (exu_idu_rf_bju_wb_preg == 6'd32) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[33] = (exu_idu_rf_bju_wb_preg == 6'd33) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[34] = (exu_idu_rf_bju_wb_preg == 6'd34) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[35] = (exu_idu_rf_bju_wb_preg == 6'd35) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[36] = (exu_idu_rf_bju_wb_preg == 6'd36) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[37] = (exu_idu_rf_bju_wb_preg == 6'd37) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[38] = (exu_idu_rf_bju_wb_preg == 6'd38) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[39] = (exu_idu_rf_bju_wb_preg == 6'd39) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[40] = (exu_idu_rf_bju_wb_preg == 6'd40) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[41] = (exu_idu_rf_bju_wb_preg == 6'd41) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[42] = (exu_idu_rf_bju_wb_preg == 6'd42) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[43] = (exu_idu_rf_bju_wb_preg == 6'd43) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[44] = (exu_idu_rf_bju_wb_preg == 6'd44) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[45] = (exu_idu_rf_bju_wb_preg == 6'd45) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[46] = (exu_idu_rf_bju_wb_preg == 6'd46) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[47] = (exu_idu_rf_bju_wb_preg == 6'd47) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[48] = (exu_idu_rf_bju_wb_preg == 6'd48) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[49] = (exu_idu_rf_bju_wb_preg == 6'd49) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[50] = (exu_idu_rf_bju_wb_preg == 6'd50) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[51] = (exu_idu_rf_bju_wb_preg == 6'd51) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[52] = (exu_idu_rf_bju_wb_preg == 6'd52) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[53] = (exu_idu_rf_bju_wb_preg == 6'd53) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[54] = (exu_idu_rf_bju_wb_preg == 6'd54) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[55] = (exu_idu_rf_bju_wb_preg == 6'd55) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[56] = (exu_idu_rf_bju_wb_preg == 6'd56) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[57] = (exu_idu_rf_bju_wb_preg == 6'd57) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[58] = (exu_idu_rf_bju_wb_preg == 6'd58) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[59] = (exu_idu_rf_bju_wb_preg == 6'd59) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[60] = (exu_idu_rf_bju_wb_preg == 6'd60) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[61] = (exu_idu_rf_bju_wb_preg == 6'd61) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[62] = (exu_idu_rf_bju_wb_preg == 6'd62) & exu_idu_rf_bju_wb_vld;
    assign bju_wb_en[63] = (exu_idu_rf_bju_wb_preg == 6'd63) & exu_idu_rf_bju_wb_vld;

    assign lsu_wb_en[0]  = (exu_idu_rf_lsu_wb_preg == 6'd0 ) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[1]  = (exu_idu_rf_lsu_wb_preg == 6'd1 ) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[2]  = (exu_idu_rf_lsu_wb_preg == 6'd2 ) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[3]  = (exu_idu_rf_lsu_wb_preg == 6'd3 ) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[4]  = (exu_idu_rf_lsu_wb_preg == 6'd4 ) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[5]  = (exu_idu_rf_lsu_wb_preg == 6'd5 ) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[6]  = (exu_idu_rf_lsu_wb_preg == 6'd6 ) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[7]  = (exu_idu_rf_lsu_wb_preg == 6'd7 ) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[8]  = (exu_idu_rf_lsu_wb_preg == 6'd8 ) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[9]  = (exu_idu_rf_lsu_wb_preg == 6'd9 ) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[10] = (exu_idu_rf_lsu_wb_preg == 6'd10) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[11] = (exu_idu_rf_lsu_wb_preg == 6'd11) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[12] = (exu_idu_rf_lsu_wb_preg == 6'd12) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[13] = (exu_idu_rf_lsu_wb_preg == 6'd13) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[14] = (exu_idu_rf_lsu_wb_preg == 6'd14) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[15] = (exu_idu_rf_lsu_wb_preg == 6'd15) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[16] = (exu_idu_rf_lsu_wb_preg == 6'd16) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[17] = (exu_idu_rf_lsu_wb_preg == 6'd17) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[18] = (exu_idu_rf_lsu_wb_preg == 6'd18) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[19] = (exu_idu_rf_lsu_wb_preg == 6'd19) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[20] = (exu_idu_rf_lsu_wb_preg == 6'd20) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[21] = (exu_idu_rf_lsu_wb_preg == 6'd21) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[22] = (exu_idu_rf_lsu_wb_preg == 6'd22) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[23] = (exu_idu_rf_lsu_wb_preg == 6'd23) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[24] = (exu_idu_rf_lsu_wb_preg == 6'd24) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[25] = (exu_idu_rf_lsu_wb_preg == 6'd25) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[26] = (exu_idu_rf_lsu_wb_preg == 6'd26) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[27] = (exu_idu_rf_lsu_wb_preg == 6'd27) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[28] = (exu_idu_rf_lsu_wb_preg == 6'd28) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[29] = (exu_idu_rf_lsu_wb_preg == 6'd29) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[30] = (exu_idu_rf_lsu_wb_preg == 6'd30) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[31] = (exu_idu_rf_lsu_wb_preg == 6'd31) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[32] = (exu_idu_rf_lsu_wb_preg == 6'd32) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[33] = (exu_idu_rf_lsu_wb_preg == 6'd33) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[34] = (exu_idu_rf_lsu_wb_preg == 6'd34) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[35] = (exu_idu_rf_lsu_wb_preg == 6'd35) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[36] = (exu_idu_rf_lsu_wb_preg == 6'd36) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[37] = (exu_idu_rf_lsu_wb_preg == 6'd37) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[38] = (exu_idu_rf_lsu_wb_preg == 6'd38) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[39] = (exu_idu_rf_lsu_wb_preg == 6'd39) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[40] = (exu_idu_rf_lsu_wb_preg == 6'd40) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[41] = (exu_idu_rf_lsu_wb_preg == 6'd41) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[42] = (exu_idu_rf_lsu_wb_preg == 6'd42) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[43] = (exu_idu_rf_lsu_wb_preg == 6'd43) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[44] = (exu_idu_rf_lsu_wb_preg == 6'd44) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[45] = (exu_idu_rf_lsu_wb_preg == 6'd45) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[46] = (exu_idu_rf_lsu_wb_preg == 6'd46) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[47] = (exu_idu_rf_lsu_wb_preg == 6'd47) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[48] = (exu_idu_rf_lsu_wb_preg == 6'd48) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[49] = (exu_idu_rf_lsu_wb_preg == 6'd49) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[50] = (exu_idu_rf_lsu_wb_preg == 6'd50) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[51] = (exu_idu_rf_lsu_wb_preg == 6'd51) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[52] = (exu_idu_rf_lsu_wb_preg == 6'd52) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[53] = (exu_idu_rf_lsu_wb_preg == 6'd53) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[54] = (exu_idu_rf_lsu_wb_preg == 6'd54) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[55] = (exu_idu_rf_lsu_wb_preg == 6'd55) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[56] = (exu_idu_rf_lsu_wb_preg == 6'd56) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[57] = (exu_idu_rf_lsu_wb_preg == 6'd57) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[58] = (exu_idu_rf_lsu_wb_preg == 6'd58) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[59] = (exu_idu_rf_lsu_wb_preg == 6'd59) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[60] = (exu_idu_rf_lsu_wb_preg == 6'd60) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[61] = (exu_idu_rf_lsu_wb_preg == 6'd61) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[62] = (exu_idu_rf_lsu_wb_preg == 6'd62) & exu_idu_rf_lsu_wb_vld;
    assign lsu_wb_en[63] = (exu_idu_rf_lsu_wb_preg == 6'd63) & exu_idu_rf_lsu_wb_vld;

    assign write_en = alu_wb_en | mxu_wb_en | div_wb_en | bju_wb_en | lsu_wb_en;
    assign write_data0  = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[0]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[0]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[0]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[0]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[0]}});
    assign write_data1  = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[1]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[1]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[1]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[1]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[1]}});
    assign write_data2  = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[2]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[2]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[2]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[2]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[2]}});
    assign write_data3  = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[3]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[3]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[3]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[3]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[3]}});
    assign write_data4  = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[4]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[4]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[4]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[4]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[4]}});
    assign write_data5  = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[5]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[5]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[5]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[5]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[5]}});
    assign write_data6  = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[6]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[6]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[6]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[6]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[6]}});
    assign write_data7  = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[7]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[7]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[7]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[7]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[7]}});
    assign write_data8  = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[8]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[8]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[8]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[8]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[8]}});
    assign write_data9  = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[9]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[9]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[9]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[9]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[9]}});
    assign write_data10 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[10]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[10]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[10]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[10]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[10]}});
    assign write_data11 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[11]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[11]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[11]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[11]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[11]}});
    assign write_data12 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[12]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[12]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[12]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[12]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[12]}});
    assign write_data13 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[13]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[13]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[13]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[13]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[13]}});
    assign write_data14 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[14]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[14]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[14]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[14]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[14]}});
    assign write_data15 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[15]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[15]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[15]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[15]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[15]}});
    assign write_data16 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[16]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[16]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[16]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[16]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[16]}});
    assign write_data17 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[17]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[17]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[17]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[17]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[17]}});
    assign write_data18 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[18]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[18]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[18]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[18]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[18]}});
    assign write_data19 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[19]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[19]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[19]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[19]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[19]}});
    assign write_data20 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[20]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[20]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[20]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[20]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[20]}});
    assign write_data21 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[21]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[21]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[21]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[21]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[21]}});
    assign write_data22 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[22]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[22]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[22]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[22]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[22]}});
    assign write_data23 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[23]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[23]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[23]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[23]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[23]}});
    assign write_data24 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[24]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[24]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[24]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[24]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[24]}});
    assign write_data25 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[25]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[25]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[25]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[25]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[25]}});
    assign write_data26 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[26]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[26]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[26]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[26]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[26]}});
    assign write_data27 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[27]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[27]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[27]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[27]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[27]}});
    assign write_data28 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[28]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[28]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[28]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[28]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[28]}});
    assign write_data29 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[29]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[29]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[29]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[29]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[29]}});
    assign write_data30 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[30]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[30]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[30]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[30]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[30]}});
    assign write_data31 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[31]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[31]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[31]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[31]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[31]}});
    assign write_data32 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[32]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[32]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[32]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[32]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[32]}});
    assign write_data33 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[33]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[33]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[33]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[33]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[33]}});
    assign write_data34 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[34]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[34]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[34]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[34]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[34]}});
    assign write_data35 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[35]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[35]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[35]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[35]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[35]}});
    assign write_data36 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[36]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[36]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[36]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[36]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[36]}});
    assign write_data37 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[37]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[37]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[37]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[37]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[37]}});
    assign write_data38 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[38]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[38]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[38]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[38]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[38]}});
    assign write_data39 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[39]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[39]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[39]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[39]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[39]}});
    assign write_data40 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[40]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[40]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[40]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[40]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[40]}});
    assign write_data41 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[41]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[41]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[41]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[41]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[41]}});
    assign write_data42 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[42]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[42]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[42]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[42]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[42]}});
    assign write_data43 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[43]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[43]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[43]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[43]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[43]}});
    assign write_data44 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[44]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[44]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[44]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[44]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[44]}});
    assign write_data45 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[45]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[45]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[45]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[45]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[45]}});
    assign write_data46 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[46]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[46]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[46]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[46]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[46]}});
    assign write_data47 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[47]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[47]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[47]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[47]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[47]}});
    assign write_data48 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[48]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[48]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[48]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[48]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[48]}});
    assign write_data49 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[49]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[49]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[49]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[49]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[49]}});
    assign write_data50 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[50]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[50]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[50]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[50]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[50]}});
    assign write_data51 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[51]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[51]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[51]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[51]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[51]}});
    assign write_data52 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[52]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[52]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[52]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[52]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[52]}});
    assign write_data53 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[53]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[53]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[53]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[53]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[53]}});
    assign write_data54 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[54]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[54]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[54]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[54]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[54]}});
    assign write_data55 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[55]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[55]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[55]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[55]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[55]}});
    assign write_data56 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[56]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[56]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[56]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[56]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[56]}});
    assign write_data57 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[57]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[57]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[57]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[57]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[57]}});
    assign write_data58 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[58]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[58]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[58]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[58]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[58]}});
    assign write_data59 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[59]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[59]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[59]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[59]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[59]}});
    assign write_data60 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[60]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[60]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[60]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[60]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[60]}});
    assign write_data61 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[61]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[61]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[61]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[61]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[61]}});
    assign write_data62 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[62]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[62]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[62]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[62]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[62]}});
    assign write_data63 = (exu_idu_rf_alu_wb_data & {64{alu_wb_en[63]}})
                        | (exu_idu_rf_mxu_wb_data & {64{mxu_wb_en[63]}})
                        | (exu_idu_rf_div_wb_data & {64{div_wb_en[63]}})
                        | (exu_idu_rf_bju_wb_data & {64{bju_wb_en[63]}})
                        | (exu_idu_rf_lsu_wb_data & {64{lsu_wb_en[63]}});
endmodule
